module foo;
endmodule

module bar;
endmodule
