module my_module();
  parameter p = q;
  parameter q = p;
endmodule
