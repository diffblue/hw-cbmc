module main;

  // reduction operators only take integral types
  wire x = &1.1;

endmodule
