module top2;
endmodule 
