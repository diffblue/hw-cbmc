module main;

  // IEEE 1800-2017 6.16
  string xyz;
  string my_string = xyz;

endmodule
