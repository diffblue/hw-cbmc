// no content

