package some_package;
  // 1800 2017 3.14.2.2
  timeunit 100ps / 10fs;
  timeprecision 10fs;
endpackage

module main;
endmodule
