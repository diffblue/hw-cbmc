module main;

  property P1;
    1
  endproperty

  assert property (P1 and P1);

endmodule
