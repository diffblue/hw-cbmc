interface myInterface;
endinterface

module main;
endmodule
