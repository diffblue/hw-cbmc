module moduleA;
endmodule

module moduleB;
endmodule
