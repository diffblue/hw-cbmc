module main(input i);

  // 1800 2017 6.20.6
  const bit my_true2 = 1;
  const var my_true3 = 1;

  // the value on the RHS does _not_ need to be constant
  const logic my_true4 = i;

endmodule
