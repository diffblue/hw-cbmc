class myClass;
endclass

module main;
  myClass x = new;
endmodule
