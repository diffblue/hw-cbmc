module main;
  wire [7:0] some_wire;
  assign some_wire[7:0] = 0;
endmodule
