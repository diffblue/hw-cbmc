module main;

  some_module_that_does_not_exist my_instance();

endmodule
