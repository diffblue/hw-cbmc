interface myInterface;
endinterface

module main;
  myInterface some_interface;
endmodule
