module top;
endmodule 

module sub;
  module nested;
  endmodule
endmodule 
