module main;
  const bit my_true2 = 1;
  const var my_true3 = 1;
  const logic my_true4 = 1;
endmodule
