module main(input clk);

  p0: assert property (0);

endmodule
