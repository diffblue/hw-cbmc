module main;
  // 'logic' is a SystemVerilog keyword
  logic some_logic;
  initial some_logic = 1;
endmodule
