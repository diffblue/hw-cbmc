module main;

  typedef struct {int a, b;} S;
  var S x = '{b:1}; // forgot a

endmodule
