module `SOME_NAME();

endmodule
