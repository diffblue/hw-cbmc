module test(some syntax error); // no newline