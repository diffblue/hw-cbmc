module main(input clk);

  p0: assert property (s_eventually 0);

endmodule
