module main;

  // % only takes integral types
  wire x = 1.1 % 1.2;

endmodule
