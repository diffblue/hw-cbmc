module main;

  wire x;

  // x is not a constant
  parameter p = x;

endmodule
