module main();

   // IEEE 1800-2017 A.2.2.1
   reg shortreal some_shortreal;
   reg real some_real;
   reg realtime some_realtime;

endmodule
