module top;
  // error: wires must have a four-valued data type
  wire bit some_wire;
endmodule
