module main;

  byte queue_of_bytes[$];
  string queue_of_strings[$:10] = { "foobar" };

endmodule
