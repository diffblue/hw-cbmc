module main;

  p0: assert final (0);

endmodule
