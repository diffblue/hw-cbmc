module main;

  always assert p0: 1 == 2;

endmodule
