module main;

  p0: assert final (real'(-1) == -1.0);

endmodule
