module main;

  parameter Q = $signed(123);

endmodule
