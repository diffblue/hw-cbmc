module main;

  // 1800-2017 6.12.1
  reg [7:0] vector;
  wire x = vector[real'(1.5)];

endmodule
