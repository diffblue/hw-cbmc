// output ports must not have a default value
module M(output [31:0] o = 4567);

endmodule
