module main;
  initial p0: assert (0);
  initial p1: assert (1);
endmodule
