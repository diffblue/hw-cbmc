module main;
  // some_var must not be redeclared
  wire [31:0] some_var;
  wire [31:0] some_var;
endmodule
