module main(input [7:0] data);

  always @(posedge data);

endmodule
