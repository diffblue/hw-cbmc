module main;

  typedef struct {int a, b;} S;
  var S x = '{b:1, something_else:0};

endmodule
