module main;

  // 1800-2017 6.12.1
  real some_real;
  wire x = some_real[0];

endmodule
