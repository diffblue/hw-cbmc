module main;

  typedef enum { E0 = 123 } my_enumt;

  assert final (E0 == 123);

endmodule
