module main;

  assert final (4'b1111 << 1 === 5'b11110);
  assert final (1 << 6 === 64);

endmodule
