module top1;
endmodule 
