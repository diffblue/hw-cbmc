module main;

  p0: assert final ('sb1 == -1);
  p1: assert final ('sb11 == -1);
  p2: assert final (4'sb111 == 7);

endmodule
