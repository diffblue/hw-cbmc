package my_package;
  typedef int some_type;
endpackage
