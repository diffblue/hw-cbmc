class myClass;
  parameter my_parameter = 123;
endclass

module main;
endmodule
