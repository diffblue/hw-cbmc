module main;

  real data;

  always @(posedge data);

endmodule
