module main(input input1);

  wire some_wire = input1;

endmodule
