module main;

  p0: assert final (real'(1'b1) == 1);

endmodule
