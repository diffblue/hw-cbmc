module main;
  assert final (0);
endmodule
