module main;

  // operand must be integral
  wire x = {<<{1.1}};

endmodule
