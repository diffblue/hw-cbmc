module main;

  // Packed arrays can be made of single bit data types
  // or other packed types.
  typedef real my_real;
  my_real [7:0] my_array;

endmodule

