module main;

  localparam x=100;

  always assert property1: x==100;

endmodule
