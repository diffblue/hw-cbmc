module main;

  function [31:0] clog2;
  input [63:0]                   value;
  reg [63:0]                     tmp;
  begin
    tmp = value - 1;
    for (clog2 = 0; tmp>0 ; clog2 = clog2 + 32'h1)
     tmp = tmp >> 1;
    end
  endfunction // clog2

  wire [clog2(16):1] x='hff; // 4 bits
  
  always assert test1: x=='b1111;

endmodule
