module main;

  reg [31:0] x;
  wire clk;

  initial expect (x==0);

endmodule
