module main;

  initial some_undeclared_task();

endmodule
