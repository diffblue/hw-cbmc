module main(x);
  // cannot declare both as input and output
  input [31:0] x;
  output [31:0] x;
endmodule
