module main();

   // IEEE 1800-2017 A.2.1.3
   var real some_real;
   var [31:0] some_word = 5;
   var signed [31:0] something_signed;
   var bit some_array[100:0];

endmodule
