module visbakery (i2,i4,i6,i8,i10,i12,i14,p0);

input i2,i4,i6,i8,i10,i12,i14;

output p0;

wire a276,a350,a414,a462,a562,a656,a884,a958,a1022,a1070,a1170,a1264,a1284,a1356,a1406,
a1426,a1454,a1482,a1518,c1,a66,a68,a70,a72,a74,a76,a78,a80,a82,a84,
a86,a88,a90,a92,a94,a96,a98,a100,a102,a104,a106,a108,a110,a112,a114,
a116,a118,a120,a122,a124,a126,a128,a130,a132,a134,a136,a138,a140,a142,a144,
a146,a148,a150,a152,a154,a156,a158,a160,a162,a164,a166,a168,a170,a172,a174,
a176,a178,a180,a182,a184,a186,a188,a190,a192,a194,a196,a198,a200,a202,a204,
a206,a208,a210,a212,a214,a216,a218,a220,a222,a224,a226,a228,a230,a232,a234,
a236,a238,a240,a242,a244,a246,a248,a250,a252,a254,a256,a258,a260,a262,a264,
a266,a268,a270,a272,a274,a278,a280,a282,a284,a286,a288,a290,a292,a294,a296,
a298,a300,a302,a304,a306,a308,a310,a312,a314,a316,a318,a320,a322,a324,a326,
a328,a330,a332,a334,a336,a338,a340,a342,a344,a346,a348,a352,a354,a356,a358,
a360,a362,a364,a366,a368,a370,a372,a374,a376,a378,a380,a382,a384,a386,a388,
a390,a392,a394,a396,a398,a400,a402,a404,a406,a408,a410,a412,a416,a418,a420,
a422,a424,a426,a428,a430,a432,a434,a436,a438,a440,a442,a444,a446,a448,a450,
a452,a454,a456,a458,a460,a464,a466,a468,a470,a472,a474,a476,a478,a480,a482,
a484,a486,a488,a490,a492,a494,a496,a498,a500,a502,a504,a506,a508,a510,a512,
a514,a516,a518,a520,a522,a524,a526,a528,a530,a532,a534,a536,a538,a540,a542,
a544,a546,a548,a550,a552,a554,a556,a558,a560,a564,a566,a568,a570,a572,a574,
a576,a578,a580,a582,a584,a586,a588,a590,a592,a594,a596,a598,a600,a602,a604,
a606,a608,a610,a612,a614,a616,a618,a620,a622,a624,a626,a628,a630,a632,a634,
a636,a638,a640,a642,a644,a646,a648,a650,a652,a654,a658,a660,a662,a664,a666,
a668,a670,a672,a674,a676,a678,a680,a682,a684,a686,a688,a690,a692,a694,a696,
a698,a700,a702,a704,a706,a708,a710,a712,a714,a716,a718,a720,a722,a724,a726,
a728,a730,a732,a734,a736,a738,a740,a742,a744,a746,a748,a750,a752,a754,a756,
a758,a760,a762,a764,a766,a768,a770,a772,a774,a776,a778,a780,a782,a784,a786,
a788,a790,a792,a794,a796,a798,a800,a802,a804,a806,a808,a810,a812,a814,a816,
a818,a820,a822,a824,a826,a828,a830,a832,a834,a836,a838,a840,a842,a844,a846,
a848,a850,a852,a854,a856,a858,a860,a862,a864,a866,a868,a870,a872,a874,a876,
a878,a880,a882,a886,a888,a890,a892,a894,a896,a898,a900,a902,a904,a906,a908,
a910,a912,a914,a916,a918,a920,a922,a924,a926,a928,a930,a932,a934,a936,a938,
a940,a942,a944,a946,a948,a950,a952,a954,a956,a960,a962,a964,a966,a968,a970,
a972,a974,a976,a978,a980,a982,a984,a986,a988,a990,a992,a994,a996,a998,a1000,
a1002,a1004,a1006,a1008,a1010,a1012,a1014,a1016,a1018,a1020,a1024,a1026,a1028,a1030,a1032,
a1034,a1036,a1038,a1040,a1042,a1044,a1046,a1048,a1050,a1052,a1054,a1056,a1058,a1060,a1062,
a1064,a1066,a1068,a1072,a1074,a1076,a1078,a1080,a1082,a1084,a1086,a1088,a1090,a1092,a1094,
a1096,a1098,a1100,a1102,a1104,a1106,a1108,a1110,a1112,a1114,a1116,a1118,a1120,a1122,a1124,
a1126,a1128,a1130,a1132,a1134,a1136,a1138,a1140,a1142,a1144,a1146,a1148,a1150,a1152,a1154,
a1156,a1158,a1160,a1162,a1164,a1166,a1168,a1172,a1174,a1176,a1178,a1180,a1182,a1184,a1186,
a1188,a1190,a1192,a1194,a1196,a1198,a1200,a1202,a1204,a1206,a1208,a1210,a1212,a1214,a1216,
a1218,a1220,a1222,a1224,a1226,a1228,a1230,a1232,a1234,a1236,a1238,a1240,a1242,a1244,a1246,
a1248,a1250,a1252,a1254,a1256,a1258,a1260,a1262,a1266,a1268,a1270,a1272,a1274,a1276,a1278,
a1280,a1282,a1286,a1288,a1290,a1292,a1294,a1296,a1298,a1300,a1302,a1304,a1306,a1308,a1310,
a1312,a1314,a1316,a1318,a1320,a1322,a1324,a1326,a1328,a1330,a1332,a1334,a1336,a1338,a1340,
a1342,a1344,a1346,a1348,a1350,a1352,a1354,a1358,a1360,a1362,a1364,a1366,a1368,a1370,a1372,
a1374,a1376,a1378,a1380,a1382,a1384,a1386,a1388,a1390,a1392,a1394,a1396,a1398,a1400,a1402,
a1404,a1408,a1410,a1412,a1414,a1416,a1418,a1420,a1422,a1424,a1428,a1430,a1432,a1434,a1436,
a1438,a1440,a1442,a1444,a1446,a1448,a1450,a1452,a1456,a1458,a1460,a1462,a1464,a1466,a1468,
a1470,a1472,a1474,a1476,a1478,a1480,a1484,a1486,a1488,a1490,a1492,a1494,a1496,a1498,a1500,
a1502,a1504,a1506,a1508,a1510,a1512,a1514,a1516,a1520,a1522,a1524,a1526,a1528,a1530,a1532,
a1534,p0;

reg l16,l18,l20,l22,l24,l26,l28,l30,l32,l34,l36,l38,l40,l42,l44,
l46,l48,l50,l52,l54,l56,l58,l60,l62,l64;

initial
begin
   l16 = 0;
   l18 = 0;
   l20 = 0;
   l22 = 0;
   l24 = 0;
   l26 = 0;
   l28 = 0;
   l30 = 0;
   l32 = 0;
   l34 = 0;
   l36 = 0;
   l38 = 0;
   l40 = 0;
   l42 = 0;
   l44 = 0;
   l46 = 0;
   l48 = 0;
   l50 = 0;
   l52 = 0;
   l54 = 0;
   l56 = 0;
   l58 = 0;
   l60 = 0;
   l62 = 0;
   l64 = 0;
end

always @(posedge i2)
   l16 <= i2;

always @(posedge i8)
   l18 <= i8;

always @(posedge i10)
   l20 <= i10;

always @(posedge a276)
   l22 <= a276;

always @(posedge a350)
   l24 <= a350;

always @(posedge a414)
   l26 <= a414;

always @(posedge a462)
   l28 <= a462;

always @(posedge a562)
   l30 <= a562;

always @(posedge a656)
   l32 <= a656;

always @(posedge a884)
   l34 <= a884;

always @(posedge a958)
   l36 <= a958;

always @(posedge a1022)
   l38 <= a1022;

always @(posedge a1070)
   l40 <= a1070;

always @(posedge a1170)
   l42 <= a1170;

always @(posedge a1264)
   l44 <= a1264;

always @(posedge i12)
   l46 <= i12;

always @(posedge i14)
   l48 <= i14;

always @(posedge a1284)
   l50 <= a1284;

always @(posedge a1356)
   l52 <= a1356;

always @(posedge a1406)
   l54 <= a1406;

always @(posedge a1426)
   l56 <= a1426;

always @(posedge a1454)
   l58 <= a1454;

always @(posedge a1482)
   l60 <= a1482;

always @(posedge a1518)
   l62 <= a1518;

always @(posedge c1)
   l64 <= c1;


assign a276 = a274 & l64;
assign a350 = a348 & l64;
assign a414 = a412 & l64;
assign a462 = a460 & l64;
assign a562 = a560 & l64;
assign a656 = a654 & l64;
assign a884 = a882 & l64;
assign a958 = a956 & l64;
assign a1022 = a1020 & l64;
assign a1070 = a1068 & l64;
assign a1170 = a1168 & l64;
assign a1264 = a1262 & l64;
assign a1284 = a1282 & l64;
assign a1356 = a1354 & l64;
assign a1406 = a1404 & l64;
assign a1426 = a1424 & l64;
assign a1454 = a1452 & l64;
assign a1482 = a1480 & l64;
assign a1518 = ~a1516 & ~a1498;
assign c1 = 1;
assign a66 = ~l22 & ~l16;
assign a68 = ~l28 & ~l26;
assign a70 = a68 & ~l24;
assign a72 = a70 & ~l22;
assign a74 = a68 & l24;
assign a76 = a74 & ~l22;
assign a78 = ~l28 & l26;
assign a80 = a78 & ~l24;
assign a82 = a80 & ~l22;
assign a84 = a78 & l24;
assign a86 = a84 & ~l22;
assign a88 = l28 & ~l26;
assign a90 = a88 & ~l24;
assign a92 = a90 & ~l22;
assign a94 = ~l32 & ~l30;
assign a96 = ~a94 & ~l50;
assign a98 = a96 & l56;
assign a100 = ~a94 & l50;
assign a102 = ~a100 & ~l56;
assign a104 = ~a102 & ~a98;
assign a106 = a88 & l24;
assign a108 = a106 & ~l22;
assign a110 = ~a94 & ~l58;
assign a112 = a110 & l52;
assign a114 = ~a94 & l58;
assign a116 = ~a114 & ~l52;
assign a118 = ~a116 & ~a112;
assign a120 = ~a94 & ~l60;
assign a122 = a120 & l54;
assign a124 = ~a94 & l60;
assign a126 = ~a124 & ~l54;
assign a128 = ~a126 & ~a122;
assign a130 = ~a128 & ~a118;
assign a132 = ~a118 & l52;
assign a134 = a132 & l54;
assign a136 = ~a134 & a128;
assign a138 = ~a132 & ~l54;
assign a140 = a138 & ~a128;
assign a142 = ~a140 & ~a136;
assign a144 = ~a118 & ~l52;
assign a146 = a118 & l52;
assign a148 = ~a146 & ~a144;
assign a150 = ~a132 & l54;
assign a152 = a132 & ~l54;
assign a154 = ~a152 & ~a150;
assign a156 = a154 & ~a128;
assign a158 = ~a154 & a128;
assign a160 = ~a158 & ~a156;
assign a162 = ~a160 & ~a148;
assign a164 = ~a162 & a142;
assign a166 = a164 & ~a130;
assign a168 = a106 & l22;
assign a170 = l28 & l26;
assign a172 = a170 & ~l24;
assign a174 = a172 & ~l22;
assign a176 = a172 & l22;
assign a178 = a170 & l24;
assign a180 = a178 & ~l22;
assign a182 = ~l22 & ~i4;
assign a184 = ~a178 & l22;
assign a186 = ~a184 & i4;
assign a188 = ~a186 & ~a182;
assign a190 = ~a188 & ~a180;
assign a192 = a190 & ~a176;
assign a194 = a192 & ~i4;
assign a196 = ~a190 & ~a176;
assign a198 = ~a196 & i4;
assign a200 = ~a198 & ~a194;
assign a202 = a200 & ~a174;
assign a204 = ~a202 & ~a168;
assign a206 = a204 & a166;
assign a208 = a202 & ~a168;
assign a210 = ~a208 & ~a166;
assign a212 = ~a210 & ~a206;
assign a214 = ~a212 & ~a108;
assign a216 = a214 & ~a104;
assign a218 = a212 & ~a108;
assign a220 = ~a218 & a104;
assign a222 = ~a220 & ~a216;
assign a224 = ~a222 & ~a92;
assign a226 = a224 & l32;
assign a228 = a222 & ~a92;
assign a230 = ~a228 & ~l32;
assign a232 = ~a230 & ~a226;
assign a234 = a232 & ~a86;
assign a236 = a234 & ~a82;
assign a238 = a236 & ~a76;
assign a240 = a238 & ~a72;
assign a242 = a240 & a66;
assign a244 = l22 & ~l16;
assign a246 = ~a244 & ~a240;
assign a248 = ~a246 & ~a242;
assign a250 = ~a178 & ~a176;
assign a252 = a250 & ~a174;
assign a254 = a252 & ~a168;
assign a256 = a254 & ~a108;
assign a258 = a256 & ~a92;
assign a260 = a258 & ~a86;
assign a262 = a260 & ~a82;
assign a264 = a262 & ~a76;
assign a266 = a264 & ~a72;
assign a268 = ~a266 & l16;
assign a270 = a268 & ~a248;
assign a272 = ~a268 & ~l22;
assign a274 = ~a272 & ~a270;
assign a278 = ~l24 & ~l16;
assign a280 = a178 & l22;
assign a282 = ~a280 & ~l24;
assign a284 = a282 & ~i4;
assign a286 = ~a280 & l24;
assign a288 = ~a286 & i4;
assign a290 = ~a288 & ~a284;
assign a292 = ~a290 & ~a180;
assign a294 = a292 & ~a176;
assign a296 = a294 & i4;
assign a298 = ~a292 & ~a176;
assign a300 = ~a298 & ~i4;
assign a302 = ~a300 & ~a296;
assign a304 = a302 & ~a174;
assign a306 = ~a304 & ~a168;
assign a308 = a306 & a166;
assign a310 = a304 & ~a168;
assign a312 = ~a310 & ~a166;
assign a314 = ~a312 & ~a308;
assign a316 = ~a314 & ~a108;
assign a318 = a316 & ~a92;
assign a320 = a318 & ~l32;
assign a322 = ~a316 & ~a92;
assign a324 = ~a322 & l32;
assign a326 = ~a324 & ~a320;
assign a328 = a326 & ~a86;
assign a330 = ~a328 & ~a82;
assign a332 = ~a330 & ~a76;
assign a334 = ~a332 & ~a72;
assign a336 = ~a334 & a278;
assign a338 = l24 & ~l16;
assign a340 = ~a338 & a334;
assign a342 = ~a340 & ~a336;
assign a344 = ~a342 & a268;
assign a346 = ~a268 & ~l24;
assign a348 = ~a346 & ~a344;
assign a352 = ~l26 & ~l16;
assign a354 = ~a280 & ~l26;
assign a356 = a354 & ~i4;
assign a358 = ~a280 & l26;
assign a360 = ~a358 & i4;
assign a362 = ~a360 & ~a356;
assign a364 = ~a362 & ~a180;
assign a366 = a364 & ~a176;
assign a368 = ~a366 & ~a174;
assign a370 = ~a368 & ~a168;
assign a372 = a370 & ~a166;
assign a374 = a368 & ~a168;
assign a376 = ~a374 & a166;
assign a378 = ~a376 & ~a372;
assign a380 = a378 & ~a108;
assign a382 = ~a380 & ~a92;
assign a384 = a382 & l32;
assign a386 = a380 & ~a92;
assign a388 = ~a386 & ~l32;
assign a390 = ~a388 & ~a384;
assign a392 = a390 & ~a86;
assign a394 = ~a392 & ~a82;
assign a396 = a394 & ~a76;
assign a398 = ~a396 & ~a72;
assign a400 = a398 & a352;
assign a402 = l26 & ~l16;
assign a404 = ~a402 & ~a398;
assign a406 = ~a404 & ~a400;
assign a408 = ~a406 & a268;
assign a410 = ~a268 & ~l26;
assign a412 = ~a410 & ~a408;
assign a416 = ~l28 & ~l16;
assign a418 = ~a280 & ~l28;
assign a420 = a418 & ~i4;
assign a422 = ~a280 & l28;
assign a424 = ~a422 & i4;
assign a426 = ~a424 & ~a420;
assign a428 = ~a426 & ~a180;
assign a430 = a428 & ~a176;
assign a432 = a430 & ~a174;
assign a434 = a432 & ~a168;
assign a436 = a434 & ~a108;
assign a438 = a436 & ~a92;
assign a440 = a438 & ~a86;
assign a442 = ~a440 & ~a82;
assign a444 = a442 & ~a76;
assign a446 = a444 & ~a72;
assign a448 = a446 & a416;
assign a450 = l28 & ~l16;
assign a452 = ~a450 & ~a446;
assign a454 = ~a452 & ~a448;
assign a456 = ~a454 & a268;
assign a458 = ~a268 & ~l28;
assign a460 = ~a458 & ~a456;
assign a464 = ~l30 & ~l16;
assign a466 = ~a174 & ~l30;
assign a468 = a174 & l30;
assign a470 = ~a468 & ~a466;
assign a472 = ~a470 & ~a168;
assign a474 = a472 & l30;
assign a476 = a470 & ~a168;
assign a478 = ~a476 & ~l30;
assign a480 = ~a478 & ~a474;
assign a482 = ~a480 & ~a108;
assign a484 = a482 & l30;
assign a486 = a480 & ~a108;
assign a488 = ~a486 & ~l30;
assign a490 = ~a488 & ~a484;
assign a492 = ~a490 & ~a92;
assign a494 = a492 & l30;
assign a496 = a490 & ~a92;
assign a498 = ~a496 & ~l30;
assign a500 = ~a498 & ~a494;
assign a502 = a500 & ~a86;
assign a504 = ~a502 & ~a82;
assign a506 = a504 & l30;
assign a508 = a502 & ~a82;
assign a510 = ~a508 & ~l30;
assign a512 = ~a510 & ~a506;
assign a514 = ~a512 & ~a76;
assign a516 = a514 & l30;
assign a518 = a512 & ~a76;
assign a520 = ~a518 & ~l30;
assign a522 = ~a520 & ~a516;
assign a524 = ~a522 & ~a72;
assign a526 = a524 & l30;
assign a528 = a522 & ~a72;
assign a530 = ~a528 & ~l30;
assign a532 = ~a530 & ~a526;
assign a534 = a532 & a464;
assign a536 = l30 & ~l16;
assign a538 = ~a536 & ~a532;
assign a540 = ~a538 & ~a534;
assign a542 = a174 & ~a106;
assign a544 = a542 & ~a92;
assign a546 = ~a544 & ~a86;
assign a548 = ~a546 & ~a82;
assign a550 = a548 & ~a76;
assign a552 = a550 & ~a72;
assign a554 = a552 & l16;
assign a556 = a554 & ~a540;
assign a558 = ~a554 & ~l30;
assign a560 = ~a558 & ~a556;
assign a564 = ~l32 & ~l16;
assign a566 = l32 & l30;
assign a568 = ~a566 & ~a94;
assign a570 = ~a174 & ~l32;
assign a572 = a570 & a568;
assign a574 = ~a174 & l32;
assign a576 = ~a574 & ~a568;
assign a578 = ~a576 & ~a572;
assign a580 = ~a578 & ~a168;
assign a582 = a580 & l32;
assign a584 = a578 & ~a168;
assign a586 = ~a584 & ~l32;
assign a588 = ~a586 & ~a582;
assign a590 = ~a588 & ~a108;
assign a592 = a590 & l32;
assign a594 = a588 & ~a108;
assign a596 = ~a594 & ~l32;
assign a598 = ~a596 & ~a592;
assign a600 = ~a598 & ~a92;
assign a602 = a600 & l32;
assign a604 = a598 & ~a92;
assign a606 = ~a604 & ~l32;
assign a608 = ~a606 & ~a602;
assign a610 = a608 & ~a86;
assign a612 = ~a610 & ~a82;
assign a614 = a612 & l32;
assign a616 = a610 & ~a82;
assign a618 = ~a616 & ~l32;
assign a620 = ~a618 & ~a614;
assign a622 = ~a620 & ~a76;
assign a624 = a622 & l32;
assign a626 = a620 & ~a76;
assign a628 = ~a626 & ~l32;
assign a630 = ~a628 & ~a624;
assign a632 = ~a630 & ~a72;
assign a634 = a632 & l32;
assign a636 = a630 & ~a72;
assign a638 = ~a636 & ~l32;
assign a640 = ~a638 & ~a634;
assign a642 = a640 & a564;
assign a644 = l32 & ~l16;
assign a646 = ~a644 & ~a640;
assign a648 = ~a646 & ~a642;
assign a650 = ~a648 & a554;
assign a652 = ~a554 & ~l32;
assign a654 = ~a652 & ~a650;
assign a658 = ~l40 & ~l38;
assign a660 = a658 & ~l36;
assign a662 = a660 & ~l34;
assign a664 = a658 & l36;
assign a666 = a664 & ~l34;
assign a668 = ~l40 & l38;
assign a670 = a668 & ~l36;
assign a672 = a670 & ~l34;
assign a674 = a668 & l36;
assign a676 = a674 & ~l34;
assign a678 = l40 & ~l38;
assign a680 = a678 & ~l36;
assign a682 = a680 & ~l34;
assign a684 = ~l44 & ~l42;
assign a686 = ~a684 & ~l50;
assign a688 = a686 & l56;
assign a690 = ~a684 & l50;
assign a692 = ~a690 & ~l56;
assign a694 = ~a692 & ~a688;
assign a696 = a678 & l36;
assign a698 = a696 & ~l34;
assign a700 = ~a684 & ~l58;
assign a702 = a700 & l52;
assign a704 = ~a684 & l58;
assign a706 = ~a704 & ~l52;
assign a708 = ~a706 & ~a702;
assign a710 = ~a684 & ~l60;
assign a712 = a710 & l54;
assign a714 = ~a684 & l60;
assign a716 = ~a714 & ~l54;
assign a718 = ~a716 & ~a712;
assign a720 = ~a718 & ~a708;
assign a722 = ~a708 & l58;
assign a724 = a722 & l60;
assign a726 = ~a724 & a718;
assign a728 = ~a722 & ~l60;
assign a730 = a728 & ~a718;
assign a732 = ~a730 & ~a726;
assign a734 = ~a708 & ~l58;
assign a736 = a708 & l58;
assign a738 = ~a736 & ~a734;
assign a740 = ~a722 & l60;
assign a742 = a722 & ~l60;
assign a744 = ~a742 & ~a740;
assign a746 = a744 & ~a718;
assign a748 = ~a744 & a718;
assign a750 = ~a748 & ~a746;
assign a752 = ~a750 & ~a738;
assign a754 = ~a752 & a732;
assign a756 = a708 & ~l58;
assign a758 = ~a756 & ~a722;
assign a760 = ~a718 & l60;
assign a762 = a718 & ~l60;
assign a764 = ~a762 & ~a760;
assign a766 = a764 & a758;
assign a768 = a766 & a684;
assign a770 = ~a768 & ~a754;
assign a772 = ~a770 & ~a720;
assign a774 = a696 & l34;
assign a776 = l40 & l38;
assign a778 = a776 & ~l36;
assign a780 = a778 & ~l34;
assign a782 = a778 & l34;
assign a784 = a776 & l36;
assign a786 = a784 & ~l34;
assign a788 = ~l34 & ~i6;
assign a790 = ~a784 & l34;
assign a792 = ~a790 & i6;
assign a794 = ~a792 & ~a788;
assign a796 = ~a794 & ~a786;
assign a798 = a796 & ~a782;
assign a800 = a798 & ~i6;
assign a802 = ~a796 & ~a782;
assign a804 = ~a802 & i6;
assign a806 = ~a804 & ~a800;
assign a808 = a806 & ~a780;
assign a810 = ~a808 & ~a774;
assign a812 = a810 & a772;
assign a814 = a808 & ~a774;
assign a816 = ~a814 & ~a772;
assign a818 = ~a816 & ~a812;
assign a820 = ~a818 & ~a698;
assign a822 = a820 & ~a694;
assign a824 = a818 & ~a698;
assign a826 = ~a824 & a694;
assign a828 = ~a826 & ~a822;
assign a830 = ~a828 & ~a682;
assign a832 = a830 & l44;
assign a834 = a828 & ~a682;
assign a836 = ~a834 & ~l44;
assign a838 = ~a836 & ~a832;
assign a840 = a838 & ~a676;
assign a842 = a840 & ~a672;
assign a844 = a842 & ~a666;
assign a846 = a844 & ~a662;
assign a848 = ~l34 & l16;
assign a850 = a848 & a846;
assign a852 = l34 & l16;
assign a854 = ~a852 & ~a846;
assign a856 = ~a854 & ~a850;
assign a858 = ~a784 & ~a782;
assign a860 = a858 & ~a780;
assign a862 = a860 & ~a774;
assign a864 = a862 & ~a698;
assign a866 = a864 & ~a682;
assign a868 = a866 & ~a676;
assign a870 = a868 & ~a672;
assign a872 = a870 & ~a666;
assign a874 = a872 & ~a662;
assign a876 = ~a874 & ~l16;
assign a878 = a876 & ~a856;
assign a880 = ~a876 & ~l34;
assign a882 = ~a880 & ~a878;
assign a886 = a784 & l34;
assign a888 = ~a886 & ~l36;
assign a890 = a888 & ~i6;
assign a892 = ~a886 & l36;
assign a894 = ~a892 & i6;
assign a896 = ~a894 & ~a890;
assign a898 = ~a896 & ~a786;
assign a900 = a898 & ~a782;
assign a902 = a900 & i6;
assign a904 = ~a898 & ~a782;
assign a906 = ~a904 & ~i6;
assign a908 = ~a906 & ~a902;
assign a910 = a908 & ~a780;
assign a912 = ~a910 & ~a774;
assign a914 = a912 & a772;
assign a916 = a910 & ~a774;
assign a918 = ~a916 & ~a772;
assign a920 = ~a918 & ~a914;
assign a922 = ~a920 & ~a698;
assign a924 = a922 & ~a682;
assign a926 = a924 & ~l44;
assign a928 = ~a922 & ~a682;
assign a930 = ~a928 & l44;
assign a932 = ~a930 & ~a926;
assign a934 = a932 & ~a676;
assign a936 = ~a934 & ~a672;
assign a938 = ~a936 & ~a666;
assign a940 = ~a938 & ~a662;
assign a942 = ~l36 & l16;
assign a944 = a942 & ~a940;
assign a946 = l36 & l16;
assign a948 = ~a946 & a940;
assign a950 = ~a948 & ~a944;
assign a952 = ~a950 & a876;
assign a954 = ~a876 & ~l36;
assign a956 = ~a954 & ~a952;
assign a960 = ~a886 & ~l38;
assign a962 = a960 & ~i6;
assign a964 = ~a886 & l38;
assign a966 = ~a964 & i6;
assign a968 = ~a966 & ~a962;
assign a970 = ~a968 & ~a786;
assign a972 = a970 & ~a782;
assign a974 = ~a972 & ~a780;
assign a976 = ~a974 & ~a774;
assign a978 = a976 & ~a772;
assign a980 = a974 & ~a774;
assign a982 = ~a980 & a772;
assign a984 = ~a982 & ~a978;
assign a986 = a984 & ~a698;
assign a988 = ~a986 & ~a682;
assign a990 = a988 & l44;
assign a992 = a986 & ~a682;
assign a994 = ~a992 & ~l44;
assign a996 = ~a994 & ~a990;
assign a998 = a996 & ~a676;
assign a1000 = ~a998 & ~a672;
assign a1002 = a1000 & ~a666;
assign a1004 = ~a1002 & ~a662;
assign a1006 = ~l38 & l16;
assign a1008 = a1006 & a1004;
assign a1010 = l38 & l16;
assign a1012 = ~a1010 & ~a1004;
assign a1014 = ~a1012 & ~a1008;
assign a1016 = ~a1014 & a876;
assign a1018 = ~a876 & ~l38;
assign a1020 = ~a1018 & ~a1016;
assign a1024 = ~a886 & ~l40;
assign a1026 = a1024 & ~i6;
assign a1028 = ~a886 & l40;
assign a1030 = ~a1028 & i6;
assign a1032 = ~a1030 & ~a1026;
assign a1034 = ~a1032 & ~a786;
assign a1036 = a1034 & ~a782;
assign a1038 = a1036 & ~a780;
assign a1040 = a1038 & ~a774;
assign a1042 = a1040 & ~a698;
assign a1044 = a1042 & ~a682;
assign a1046 = a1044 & ~a676;
assign a1048 = ~a1046 & ~a672;
assign a1050 = a1048 & ~a666;
assign a1052 = a1050 & ~a662;
assign a1054 = ~l40 & l16;
assign a1056 = a1054 & a1052;
assign a1058 = l40 & l16;
assign a1060 = ~a1058 & ~a1052;
assign a1062 = ~a1060 & ~a1056;
assign a1064 = ~a1062 & a876;
assign a1066 = ~a876 & ~l40;
assign a1068 = ~a1066 & ~a1064;
assign a1072 = ~a780 & ~l42;
assign a1074 = a780 & l42;
assign a1076 = ~a1074 & ~a1072;
assign a1078 = ~a1076 & ~a774;
assign a1080 = a1078 & l42;
assign a1082 = a1076 & ~a774;
assign a1084 = ~a1082 & ~l42;
assign a1086 = ~a1084 & ~a1080;
assign a1088 = ~a1086 & ~a698;
assign a1090 = a1088 & l42;
assign a1092 = a1086 & ~a698;
assign a1094 = ~a1092 & ~l42;
assign a1096 = ~a1094 & ~a1090;
assign a1098 = ~a1096 & ~a682;
assign a1100 = a1098 & l42;
assign a1102 = a1096 & ~a682;
assign a1104 = ~a1102 & ~l42;
assign a1106 = ~a1104 & ~a1100;
assign a1108 = a1106 & ~a676;
assign a1110 = ~a1108 & ~a672;
assign a1112 = a1110 & l42;
assign a1114 = a1108 & ~a672;
assign a1116 = ~a1114 & ~l42;
assign a1118 = ~a1116 & ~a1112;
assign a1120 = ~a1118 & ~a666;
assign a1122 = a1120 & l42;
assign a1124 = a1118 & ~a666;
assign a1126 = ~a1124 & ~l42;
assign a1128 = ~a1126 & ~a1122;
assign a1130 = ~a1128 & ~a662;
assign a1132 = a1130 & l42;
assign a1134 = a1128 & ~a662;
assign a1136 = ~a1134 & ~l42;
assign a1138 = ~a1136 & ~a1132;
assign a1140 = ~l42 & l16;
assign a1142 = a1140 & a1138;
assign a1144 = l42 & l16;
assign a1146 = ~a1144 & ~a1138;
assign a1148 = ~a1146 & ~a1142;
assign a1150 = a780 & ~a696;
assign a1152 = a1150 & ~a682;
assign a1154 = ~a1152 & ~a676;
assign a1156 = ~a1154 & ~a672;
assign a1158 = a1156 & ~a666;
assign a1160 = a1158 & ~a662;
assign a1162 = a1160 & ~l16;
assign a1164 = a1162 & ~a1148;
assign a1166 = ~a1162 & ~l42;
assign a1168 = ~a1166 & ~a1164;
assign a1172 = l44 & l42;
assign a1174 = ~a1172 & ~a684;
assign a1176 = ~a780 & ~l44;
assign a1178 = a1176 & a1174;
assign a1180 = ~a780 & l44;
assign a1182 = ~a1180 & ~a1174;
assign a1184 = ~a1182 & ~a1178;
assign a1186 = ~a1184 & ~a774;
assign a1188 = a1186 & l44;
assign a1190 = a1184 & ~a774;
assign a1192 = ~a1190 & ~l44;
assign a1194 = ~a1192 & ~a1188;
assign a1196 = ~a1194 & ~a698;
assign a1198 = a1196 & l44;
assign a1200 = a1194 & ~a698;
assign a1202 = ~a1200 & ~l44;
assign a1204 = ~a1202 & ~a1198;
assign a1206 = ~a1204 & ~a682;
assign a1208 = a1206 & l44;
assign a1210 = a1204 & ~a682;
assign a1212 = ~a1210 & ~l44;
assign a1214 = ~a1212 & ~a1208;
assign a1216 = a1214 & ~a676;
assign a1218 = ~a1216 & ~a672;
assign a1220 = a1218 & l44;
assign a1222 = a1216 & ~a672;
assign a1224 = ~a1222 & ~l44;
assign a1226 = ~a1224 & ~a1220;
assign a1228 = ~a1226 & ~a666;
assign a1230 = a1228 & l44;
assign a1232 = a1226 & ~a666;
assign a1234 = ~a1232 & ~l44;
assign a1236 = ~a1234 & ~a1230;
assign a1238 = ~a1236 & ~a662;
assign a1240 = a1238 & l44;
assign a1242 = a1236 & ~a662;
assign a1244 = ~a1242 & ~l44;
assign a1246 = ~a1244 & ~a1240;
assign a1248 = ~l44 & l16;
assign a1250 = a1248 & a1246;
assign a1252 = l44 & l16;
assign a1254 = ~a1252 & ~a1246;
assign a1256 = ~a1254 & ~a1250;
assign a1258 = ~a1256 & a1162;
assign a1260 = ~a1162 & ~l44;
assign a1262 = ~a1260 & ~a1258;
assign a1266 = ~l50 & l16;
assign a1268 = ~a672 & l50;
assign a1270 = ~a1268 & ~a662;
assign a1272 = ~a1270 & a1266;
assign a1274 = l50 & l16;
assign a1276 = ~a1274 & a1270;
assign a1278 = ~a1276 & ~a1272;
assign a1280 = ~a1278 & ~l16;
assign a1282 = ~a1280 & ~a1266;
assign a1286 = ~l52 & ~l16;
assign a1288 = l58 & ~l52;
assign a1290 = a1288 & l60;
assign a1292 = ~a1290 & l54;
assign a1294 = ~a1288 & ~l60;
assign a1296 = a1294 & ~l54;
assign a1298 = ~a1296 & ~a1292;
assign a1300 = ~l58 & ~l52;
assign a1302 = l58 & l52;
assign a1304 = ~a1302 & ~a1300;
assign a1306 = a1288 & ~l60;
assign a1308 = ~a1288 & l60;
assign a1310 = ~a1308 & ~a1306;
assign a1312 = a1310 & ~l54;
assign a1314 = ~a1310 & l54;
assign a1316 = ~a1314 & ~a1312;
assign a1318 = ~a1316 & ~a1304;
assign a1320 = ~a1318 & ~a1298;
assign a1322 = ~a1320 & l58;
assign a1324 = a1322 & ~l52;
assign a1326 = ~a1320 & ~l58;
assign a1328 = ~a1326 & l52;
assign a1330 = ~a1328 & ~a1324;
assign a1332 = ~a76 & ~l52;
assign a1334 = a1332 & a1330;
assign a1336 = ~a76 & l52;
assign a1338 = ~a1336 & ~a1330;
assign a1340 = ~a1338 & ~a1334;
assign a1342 = a1340 & ~a180;
assign a1344 = a1342 & a1286;
assign a1346 = l52 & ~l16;
assign a1348 = ~a1346 & ~a1342;
assign a1350 = ~a1348 & ~a1344;
assign a1352 = ~a1350 & l16;
assign a1354 = ~a1352 & ~a1286;
assign a1358 = ~l54 & ~l16;
assign a1360 = ~l54 & ~l52;
assign a1362 = l54 & l52;
assign a1364 = ~a1362 & ~a1360;
assign a1366 = ~l60 & ~l58;
assign a1368 = l60 & l58;
assign a1370 = ~a1368 & ~a1366;
assign a1372 = ~a1370 & ~a1320;
assign a1374 = a1372 & a1364;
assign a1376 = a1370 & ~a1320;
assign a1378 = ~a1376 & ~a1364;
assign a1380 = ~a1378 & ~a1374;
assign a1382 = ~a76 & ~l54;
assign a1384 = a1382 & a1380;
assign a1386 = ~a76 & l54;
assign a1388 = ~a1386 & ~a1380;
assign a1390 = ~a1388 & ~a1384;
assign a1392 = a1390 & ~a180;
assign a1394 = a1392 & a1358;
assign a1396 = l54 & ~l16;
assign a1398 = ~a1396 & ~a1392;
assign a1400 = ~a1398 & ~a1394;
assign a1402 = ~a1400 & l16;
assign a1404 = ~a1402 & ~a1358;
assign a1408 = ~l56 & ~l16;
assign a1410 = ~a82 & l56;
assign a1412 = ~a1410 & ~a72;
assign a1414 = ~a1412 & a1408;
assign a1416 = l56 & ~l16;
assign a1418 = ~a1416 & a1412;
assign a1420 = ~a1418 & ~a1414;
assign a1422 = ~a1420 & l16;
assign a1424 = ~a1422 & ~a1408;
assign a1428 = ~l58 & l16;
assign a1430 = ~a666 & ~l58;
assign a1432 = a1430 & a1330;
assign a1434 = ~a666 & l58;
assign a1436 = ~a1434 & ~a1330;
assign a1438 = ~a1436 & ~a1432;
assign a1440 = a1438 & ~a786;
assign a1442 = a1440 & a1428;
assign a1444 = l58 & l16;
assign a1446 = ~a1444 & ~a1440;
assign a1448 = ~a1446 & ~a1442;
assign a1450 = ~a1448 & ~l16;
assign a1452 = ~a1450 & ~a1428;
assign a1456 = ~l60 & l16;
assign a1458 = ~a666 & ~l60;
assign a1460 = a1458 & a1380;
assign a1462 = ~a666 & l60;
assign a1464 = ~a1462 & ~a1380;
assign a1466 = ~a1464 & ~a1460;
assign a1468 = a1466 & ~a786;
assign a1470 = a1468 & a1456;
assign a1472 = l60 & l16;
assign a1474 = ~a1472 & ~a1468;
assign a1476 = ~a1474 & ~a1470;
assign a1478 = ~a1476 & ~l16;
assign a1480 = ~a1478 & ~a1456;
assign a1484 = ~i12 & i10;
assign a1486 = i12 & ~i10;
assign a1488 = ~a1486 & ~a1484;
assign a1490 = ~i14 & i8;
assign a1492 = i14 & ~i8;
assign a1494 = ~a1492 & ~a1490;
assign a1496 = a1494 & a1488;
assign a1498 = ~a1496 & ~l64;
assign a1500 = ~l16 & ~i12;
assign a1502 = l16 & i12;
assign a1504 = ~a1502 & ~a1500;
assign a1506 = l16 & ~i14;
assign a1508 = ~l16 & i14;
assign a1510 = ~a1508 & ~a1506;
assign a1512 = a1510 & a1504;
assign a1514 = a1512 & l62;
assign a1516 = ~a1514 & l64;
assign a1520 = ~l24 & l22;
assign a1522 = a1520 & l26;
assign a1524 = a1522 & l28;
assign a1526 = ~l36 & l34;
assign a1528 = a1526 & l38;
assign a1530 = a1528 & l40;
assign a1532 = a1530 & a1524;
assign a1534 = a1532 & l62;
assign p0 = a1534;

assert property (~p0);

endmodule
