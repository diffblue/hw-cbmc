module main;

  reg [7:0] my_array[10] = '{1, 2, 3, 4}; // too short

endmodule
