module ;// forgot the name
