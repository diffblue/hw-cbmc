module main;

  wire [31:0] x = {4{1.1}};

endmodule
