module main;

  // arithmetic shift
  assert final (-1 >>> 1 === -1);
  assert final (1 >>> 1 === 0);
  assert final (-2 >>> 1 === -1);

endmodule
