module main;

  // no synthesis semantics at all
  final $display("Final time: %d", $time);

endmodule
