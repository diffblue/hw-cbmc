module main(input [31:0] some_var);
  // some_var must not be redeclared
  input [31:0] some_var;
endmodule
