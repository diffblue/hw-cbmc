module main(; // forgot the )
