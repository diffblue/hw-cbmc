module main(input clk);

  initial p0: assert property (0);

endmodule
