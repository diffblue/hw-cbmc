module main;

  wire y = this;

endmodule
