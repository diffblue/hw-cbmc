module main // forgot the ;

byte some_var;

endmodule

