module my_module(some_port);

  // some_port is not declared as input or output

endmodule
