class myClass;
  parameter my_parameter = 123;
endclass

module main;
  myClass c = null;
endmodule
