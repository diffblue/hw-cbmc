module sm98a7multi (i2,i4,i6,i8,i10,i12,i14,i16,i18,i20,i22,i24,i26,i28,i30,
i32,i34,i36,i38,i40,i42,i44,i46,i48,i50,i52,i54,i56,i58,i60,
i62,i64,i66,i68,i70,i72,i74,i76,i78,i80,i82,i84,i86,i88,i90,
i92,i94,i96,i98,i100,i102,i104,i106,i108,i110,i112,i114,i116,i118,i120,
i122,i124,i126,i128,i130,i132,i134,i136,i138,i140,i142,i144,i146,i148,i150,
i152,i154,i156,i158,i160,i162,p0,p1,p2,p3,p4);

input i2,i4,i6,i8,i10,i12,i14,i16,i18,i20,i22,i24,i26,i28,i30,
i32,i34,i36,i38,i40,i42,i44,i46,i48,i50,i52,i54,i56,i58,i60,
i62,i64,i66,i68,i70,i72,i74,i76,i78,i80,i82,i84,i86,i88,i90,
i92,i94,i96,i98,i100,i102,i104,i106,i108,i110,i112,i114,i116,i118,i120,
i122,i124,i126,i128,i130,i132,i134,i136,i138,i140,i142,i144,i146,i148,i150,
i152,i154,i156,i158,i160,i162;

output p0,p1,p2,p3,p4;

wire na342,a344,na346,a348,a350,z0,a19472,c1,a342,a346,a352,a354,a356,a358,a360,
a362,a364,a366,a368,a370,a372,a374,a376,a378,a380,a382,a384,a386,a388,a390,
a392,a394,a396,a398,a400,a402,a404,a406,a408,a410,a412,a414,a416,a418,a420,
a422,a424,a426,a428,a430,a432,a434,a436,a438,a440,a442,a444,a446,a448,a450,
a452,a454,a456,a458,a460,a462,a464,a466,a468,a470,a472,a474,a476,a478,a480,
a482,a484,a486,a488,a490,a492,a494,a496,a498,a500,a502,a504,a506,a508,a510,
a512,a514,a516,a518,a520,a522,a524,a526,a528,a530,a532,a534,a536,a538,a540,
a542,a544,a546,a548,a550,a552,a554,a556,a558,a560,a562,a564,a566,a568,a570,
a572,a574,a576,a578,a580,a582,a584,a586,a588,a590,a592,a594,a596,a598,a600,
a602,a604,a606,a608,a610,a612,a614,a616,a618,a620,a622,a624,a626,a628,a630,
a632,a634,a636,a638,a640,a642,a644,a646,a648,a650,a652,a654,a656,a658,a660,
a662,a664,a666,a668,a670,a672,a674,a676,a678,a680,a682,a684,a686,a688,a690,
a692,a694,a696,a698,a700,a702,a704,a706,a708,a710,a712,a714,a716,a718,a720,
a722,a724,a726,a728,a730,a732,a734,a736,a738,a740,a742,a744,a746,a748,a750,
a752,a754,a756,a758,a760,a762,a764,a766,a768,a770,a772,a774,a776,a778,a780,
a782,a784,a786,a788,a790,a792,a794,a796,a798,a800,a802,a804,a806,a808,a810,
a812,a814,a816,a818,a820,a822,a824,a826,a828,a830,a832,a834,a836,a838,a840,
a842,a844,a846,a848,a850,a852,a854,a856,a858,a860,a862,a864,a866,a868,a870,
a872,a874,a876,a878,a880,a882,a884,a886,a888,a890,a892,a894,a896,a898,a900,
a902,a904,a906,a908,a910,a912,a914,a916,a918,a920,a922,a924,a926,a928,a930,
a932,a934,a936,a938,a940,a942,a944,a946,a948,a950,a952,a954,a956,a958,a960,
a962,a964,a966,a968,a970,a972,a974,a976,a978,a980,a982,a984,a986,a988,a990,
a992,a994,a996,a998,a1000,a1002,a1004,a1006,a1008,a1010,a1012,a1014,a1016,a1018,a1020,
a1022,a1024,a1026,a1028,a1030,a1032,a1034,a1036,a1038,a1040,a1042,a1044,a1046,a1048,a1050,
a1052,a1054,a1056,a1058,a1060,a1062,a1064,a1066,a1068,a1070,a1072,a1074,a1076,a1078,a1080,
a1082,a1084,a1086,a1088,a1090,a1092,a1094,a1096,a1098,a1100,a1102,a1104,a1106,a1108,a1110,
a1112,a1114,a1116,a1118,a1120,a1122,a1124,a1126,a1128,a1130,a1132,a1134,a1136,a1138,a1140,
a1142,a1144,a1146,a1148,a1150,a1152,a1154,a1156,a1158,a1160,a1162,a1164,a1166,a1168,a1170,
a1172,a1174,a1176,a1178,a1180,a1182,a1184,a1186,a1188,a1190,a1192,a1194,a1196,a1198,a1200,
a1202,a1204,a1206,a1208,a1210,a1212,a1214,a1216,a1218,a1220,a1222,a1224,a1226,a1228,a1230,
a1232,a1234,a1236,a1238,a1240,a1242,a1244,a1246,a1248,a1250,a1252,a1254,a1256,a1258,a1260,
a1262,a1264,a1266,a1268,a1270,a1272,a1274,a1276,a1278,a1280,a1282,a1284,a1286,a1288,a1290,
a1292,a1294,a1296,a1298,a1300,a1302,a1304,a1306,a1308,a1310,a1312,a1314,a1316,a1318,a1320,
a1322,a1324,a1326,a1328,a1330,a1332,a1334,a1336,a1338,a1340,a1342,a1344,a1346,a1348,a1350,
a1352,a1354,a1356,a1358,a1360,a1362,a1364,a1366,a1368,a1370,a1372,a1374,a1376,a1378,a1380,
a1382,a1384,a1386,a1388,a1390,a1392,a1394,a1396,a1398,a1400,a1402,a1404,a1406,a1408,a1410,
a1412,a1414,a1416,a1418,a1420,a1422,a1424,a1426,a1428,a1430,a1432,a1434,a1436,a1438,a1440,
a1442,a1444,a1446,a1448,a1450,a1452,a1454,a1456,a1458,a1460,a1462,a1464,a1466,a1468,a1470,
a1472,a1474,a1476,a1478,a1480,a1482,a1484,a1486,a1488,a1490,a1492,a1494,a1496,a1498,a1500,
a1502,a1504,a1506,a1508,a1510,a1512,a1514,a1516,a1518,a1520,a1522,a1524,a1526,a1528,a1530,
a1532,a1534,a1536,a1538,a1540,a1542,a1544,a1546,a1548,a1550,a1552,a1554,a1556,a1558,a1560,
a1562,a1564,a1566,a1568,a1570,a1572,a1574,a1576,a1578,a1580,a1582,a1584,a1586,a1588,a1590,
a1592,a1594,a1596,a1598,a1600,a1602,a1604,a1606,a1608,a1610,a1612,a1614,a1616,a1618,a1620,
a1622,a1624,a1626,a1628,a1630,a1632,a1634,a1636,a1638,a1640,a1642,a1644,a1646,a1648,a1650,
a1652,a1654,a1656,a1658,a1660,a1662,a1664,a1666,a1668,a1670,a1672,a1674,a1676,a1678,a1680,
a1682,a1684,a1686,a1688,a1690,a1692,a1694,a1696,a1698,a1700,a1702,a1704,a1706,a1708,a1710,
a1712,a1714,a1716,a1718,a1720,a1722,a1724,a1726,a1728,a1730,a1732,a1734,a1736,a1738,a1740,
a1742,a1744,a1746,a1748,a1750,a1752,a1754,a1756,a1758,a1760,a1762,a1764,a1766,a1768,a1770,
a1772,a1774,a1776,a1778,a1780,a1782,a1784,a1786,a1788,a1790,a1792,a1794,a1796,a1798,a1800,
a1802,a1804,a1806,a1808,a1810,a1812,a1814,a1816,a1818,a1820,a1822,a1824,a1826,a1828,a1830,
a1832,a1834,a1836,a1838,a1840,a1842,a1844,a1846,a1848,a1850,a1852,a1854,a1856,a1858,a1860,
a1862,a1864,a1866,a1868,a1870,a1872,a1874,a1876,a1878,a1880,a1882,a1884,a1886,a1888,a1890,
a1892,a1894,a1896,a1898,a1900,a1902,a1904,a1906,a1908,a1910,a1912,a1914,a1916,a1918,a1920,
a1922,a1924,a1926,a1928,a1930,a1932,a1934,a1936,a1938,a1940,a1942,a1944,a1946,a1948,a1950,
a1952,a1954,a1956,a1958,a1960,a1962,a1964,a1966,a1968,a1970,a1972,a1974,a1976,a1978,a1980,
a1982,a1984,a1986,a1988,a1990,a1992,a1994,a1996,a1998,a2000,a2002,a2004,a2006,a2008,a2010,
a2012,a2014,a2016,a2018,a2020,a2022,a2024,a2026,a2028,a2030,a2032,a2034,a2036,a2038,a2040,
a2042,a2044,a2046,a2048,a2050,a2052,a2054,a2056,a2058,a2060,a2062,a2064,a2066,a2068,a2070,
a2072,a2074,a2076,a2078,a2080,a2082,a2084,a2086,a2088,a2090,a2092,a2094,a2096,a2098,a2100,
a2102,a2104,a2106,a2108,a2110,a2112,a2114,a2116,a2118,a2120,a2122,a2124,a2126,a2128,a2130,
a2132,a2134,a2136,a2138,a2140,a2142,a2144,a2146,a2148,a2150,a2152,a2154,a2156,a2158,a2160,
a2162,a2164,a2166,a2168,a2170,a2172,a2174,a2176,a2178,a2180,a2182,a2184,a2186,a2188,a2190,
a2192,a2194,a2196,a2198,a2200,a2202,a2204,a2206,a2208,a2210,a2212,a2214,a2216,a2218,a2220,
a2222,a2224,a2226,a2228,a2230,a2232,a2234,a2236,a2238,a2240,a2242,a2244,a2246,a2248,a2250,
a2252,a2254,a2256,a2258,a2260,a2262,a2264,a2266,a2268,a2270,a2272,a2274,a2276,a2278,a2280,
a2282,a2284,a2286,a2288,a2290,a2292,a2294,a2296,a2298,a2300,a2302,a2304,a2306,a2308,a2310,
a2312,a2314,a2316,a2318,a2320,a2322,a2324,a2326,a2328,a2330,a2332,a2334,a2336,a2338,a2340,
a2342,a2344,a2346,a2348,a2350,a2352,a2354,a2356,a2358,a2360,a2362,a2364,a2366,a2368,a2370,
a2372,a2374,a2376,a2378,a2380,a2382,a2384,a2386,a2388,a2390,a2392,a2394,a2396,a2398,a2400,
a2402,a2404,a2406,a2408,a2410,a2412,a2414,a2416,a2418,a2420,a2422,a2424,a2426,a2428,a2430,
a2432,a2434,a2436,a2438,a2440,a2442,a2444,a2446,a2448,a2450,a2452,a2454,a2456,a2458,a2460,
a2462,a2464,a2466,a2468,a2470,a2472,a2474,a2476,a2478,a2480,a2482,a2484,a2486,a2488,a2490,
a2492,a2494,a2496,a2498,a2500,a2502,a2504,a2506,a2508,a2510,a2512,a2514,a2516,a2518,a2520,
a2522,a2524,a2526,a2528,a2530,a2532,a2534,a2536,a2538,a2540,a2542,a2544,a2546,a2548,a2550,
a2552,a2554,a2556,a2558,a2560,a2562,a2564,a2566,a2568,a2570,a2572,a2574,a2576,a2578,a2580,
a2582,a2584,a2586,a2588,a2590,a2592,a2594,a2596,a2598,a2600,a2602,a2604,a2606,a2608,a2610,
a2612,a2614,a2616,a2618,a2620,a2622,a2624,a2626,a2628,a2630,a2632,a2634,a2636,a2638,a2640,
a2642,a2644,a2646,a2648,a2650,a2652,a2654,a2656,a2658,a2660,a2662,a2664,a2666,a2668,a2670,
a2672,a2674,a2676,a2678,a2680,a2682,a2684,a2686,a2688,a2690,a2692,a2694,a2696,a2698,a2700,
a2702,a2704,a2706,a2708,a2710,a2712,a2714,a2716,a2718,a2720,a2722,a2724,a2726,a2728,a2730,
a2732,a2734,a2736,a2738,a2740,a2742,a2744,a2746,a2748,a2750,a2752,a2754,a2756,a2758,a2760,
a2762,a2764,a2766,a2768,a2770,a2772,a2774,a2776,a2778,a2780,a2782,a2784,a2786,a2788,a2790,
a2792,a2794,a2796,a2798,a2800,a2802,a2804,a2806,a2808,a2810,a2812,a2814,a2816,a2818,a2820,
a2822,a2824,a2826,a2828,a2830,a2832,a2834,a2836,a2838,a2840,a2842,a2844,a2846,a2848,a2850,
a2852,a2854,a2856,a2858,a2860,a2862,a2864,a2866,a2868,a2870,a2872,a2874,a2876,a2878,a2880,
a2882,a2884,a2886,a2888,a2890,a2892,a2894,a2896,a2898,a2900,a2902,a2904,a2906,a2908,a2910,
a2912,a2914,a2916,a2918,a2920,a2922,a2924,a2926,a2928,a2930,a2932,a2934,a2936,a2938,a2940,
a2942,a2944,a2946,a2948,a2950,a2952,a2954,a2956,a2958,a2960,a2962,a2964,a2966,a2968,a2970,
a2972,a2974,a2976,a2978,a2980,a2982,a2984,a2986,a2988,a2990,a2992,a2994,a2996,a2998,a3000,
a3002,a3004,a3006,a3008,a3010,a3012,a3014,a3016,a3018,a3020,a3022,a3024,a3026,a3028,a3030,
a3032,a3034,a3036,a3038,a3040,a3042,a3044,a3046,a3048,a3050,a3052,a3054,a3056,a3058,a3060,
a3062,a3064,a3066,a3068,a3070,a3072,a3074,a3076,a3078,a3080,a3082,a3084,a3086,a3088,a3090,
a3092,a3094,a3096,a3098,a3100,a3102,a3104,a3106,a3108,a3110,a3112,a3114,a3116,a3118,a3120,
a3122,a3124,a3126,a3128,a3130,a3132,a3134,a3136,a3138,a3140,a3142,a3144,a3146,a3148,a3150,
a3152,a3154,a3156,a3158,a3160,a3162,a3164,a3166,a3168,a3170,a3172,a3174,a3176,a3178,a3180,
a3182,a3184,a3186,a3188,a3190,a3192,a3194,a3196,a3198,a3200,a3202,a3204,a3206,a3208,a3210,
a3212,a3214,a3216,a3218,a3220,a3222,a3224,a3226,a3228,a3230,a3232,a3234,a3236,a3238,a3240,
a3242,a3244,a3246,a3248,a3250,a3252,a3254,a3256,a3258,a3260,a3262,a3264,a3266,a3268,a3270,
a3272,a3274,a3276,a3278,a3280,a3282,a3284,a3286,a3288,a3290,a3292,a3294,a3296,a3298,a3300,
a3302,a3304,a3306,a3308,a3310,a3312,a3314,a3316,a3318,a3320,a3322,a3324,a3326,a3328,a3330,
a3332,a3334,a3336,a3338,a3340,a3342,a3344,a3346,a3348,a3350,a3352,a3354,a3356,a3358,a3360,
a3362,a3364,a3366,a3368,a3370,a3372,a3374,a3376,a3378,a3380,a3382,a3384,a3386,a3388,a3390,
a3392,a3394,a3396,a3398,a3400,a3402,a3404,a3406,a3408,a3410,a3412,a3414,a3416,a3418,a3420,
a3422,a3424,a3426,a3428,a3430,a3432,a3434,a3436,a3438,a3440,a3442,a3444,a3446,a3448,a3450,
a3452,a3454,a3456,a3458,a3460,a3462,a3464,a3466,a3468,a3470,a3472,a3474,a3476,a3478,a3480,
a3482,a3484,a3486,a3488,a3490,a3492,a3494,a3496,a3498,a3500,a3502,a3504,a3506,a3508,a3510,
a3512,a3514,a3516,a3518,a3520,a3522,a3524,a3526,a3528,a3530,a3532,a3534,a3536,a3538,a3540,
a3542,a3544,a3546,a3548,a3550,a3552,a3554,a3556,a3558,a3560,a3562,a3564,a3566,a3568,a3570,
a3572,a3574,a3576,a3578,a3580,a3582,a3584,a3586,a3588,a3590,a3592,a3594,a3596,a3598,a3600,
a3602,a3604,a3606,a3608,a3610,a3612,a3614,a3616,a3618,a3620,a3622,a3624,a3626,a3628,a3630,
a3632,a3634,a3636,a3638,a3640,a3642,a3644,a3646,a3648,a3650,a3652,a3654,a3656,a3658,a3660,
a3662,a3664,a3666,a3668,a3670,a3672,a3674,a3676,a3678,a3680,a3682,a3684,a3686,a3688,a3690,
a3692,a3694,a3696,a3698,a3700,a3702,a3704,a3706,a3708,a3710,a3712,a3714,a3716,a3718,a3720,
a3722,a3724,a3726,a3728,a3730,a3732,a3734,a3736,a3738,a3740,a3742,a3744,a3746,a3748,a3750,
a3752,a3754,a3756,a3758,a3760,a3762,a3764,a3766,a3768,a3770,a3772,a3774,a3776,a3778,a3780,
a3782,a3784,a3786,a3788,a3790,a3792,a3794,a3796,a3798,a3800,a3802,a3804,a3806,a3808,a3810,
a3812,a3814,a3816,a3818,a3820,a3822,a3824,a3826,a3828,a3830,a3832,a3834,a3836,a3838,a3840,
a3842,a3844,a3846,a3848,a3850,a3852,a3854,a3856,a3858,a3860,a3862,a3864,a3866,a3868,a3870,
a3872,a3874,a3876,a3878,a3880,a3882,a3884,a3886,a3888,a3890,a3892,a3894,a3896,a3898,a3900,
a3902,a3904,a3906,a3908,a3910,a3912,a3914,a3916,a3918,a3920,a3922,a3924,a3926,a3928,a3930,
a3932,a3934,a3936,a3938,a3940,a3942,a3944,a3946,a3948,a3950,a3952,a3954,a3956,a3958,a3960,
a3962,a3964,a3966,a3968,a3970,a3972,a3974,a3976,a3978,a3980,a3982,a3984,a3986,a3988,a3990,
a3992,a3994,a3996,a3998,a4000,a4002,a4004,a4006,a4008,a4010,a4012,a4014,a4016,a4018,a4020,
a4022,a4024,a4026,a4028,a4030,a4032,a4034,a4036,a4038,a4040,a4042,a4044,a4046,a4048,a4050,
a4052,a4054,a4056,a4058,a4060,a4062,a4064,a4066,a4068,a4070,a4072,a4074,a4076,a4078,a4080,
a4082,a4084,a4086,a4088,a4090,a4092,a4094,a4096,a4098,a4100,a4102,a4104,a4106,a4108,a4110,
a4112,a4114,a4116,a4118,a4120,a4122,a4124,a4126,a4128,a4130,a4132,a4134,a4136,a4138,a4140,
a4142,a4144,a4146,a4148,a4150,a4152,a4154,a4156,a4158,a4160,a4162,a4164,a4166,a4168,a4170,
a4172,a4174,a4176,a4178,a4180,a4182,a4184,a4186,a4188,a4190,a4192,a4194,a4196,a4198,a4200,
a4202,a4204,a4206,a4208,a4210,a4212,a4214,a4216,a4218,a4220,a4222,a4224,a4226,a4228,a4230,
a4232,a4234,a4236,a4238,a4240,a4242,a4244,a4246,a4248,a4250,a4252,a4254,a4256,a4258,a4260,
a4262,a4264,a4266,a4268,a4270,a4272,a4274,a4276,a4278,a4280,a4282,a4284,a4286,a4288,a4290,
a4292,a4294,a4296,a4298,a4300,a4302,a4304,a4306,a4308,a4310,a4312,a4314,a4316,a4318,a4320,
a4322,a4324,a4326,a4328,a4330,a4332,a4334,a4336,a4338,a4340,a4342,a4344,a4346,a4348,a4350,
a4352,a4354,a4356,a4358,a4360,a4362,a4364,a4366,a4368,a4370,a4372,a4374,a4376,a4378,a4380,
a4382,a4384,a4386,a4388,a4390,a4392,a4394,a4396,a4398,a4400,a4402,a4404,a4406,a4408,a4410,
a4412,a4414,a4416,a4418,a4420,a4422,a4424,a4426,a4428,a4430,a4432,a4434,a4436,a4438,a4440,
a4442,a4444,a4446,a4448,a4450,a4452,a4454,a4456,a4458,a4460,a4462,a4464,a4466,a4468,a4470,
a4472,a4474,a4476,a4478,a4480,a4482,a4484,a4486,a4488,a4490,a4492,a4494,a4496,a4498,a4500,
a4502,a4504,a4506,a4508,a4510,a4512,a4514,a4516,a4518,a4520,a4522,a4524,a4526,a4528,a4530,
a4532,a4534,a4536,a4538,a4540,a4542,a4544,a4546,a4548,a4550,a4552,a4554,a4556,a4558,a4560,
a4562,a4564,a4566,a4568,a4570,a4572,a4574,a4576,a4578,a4580,a4582,a4584,a4586,a4588,a4590,
a4592,a4594,a4596,a4598,a4600,a4602,a4604,a4606,a4608,a4610,a4612,a4614,a4616,a4618,a4620,
a4622,a4624,a4626,a4628,a4630,a4632,a4634,a4636,a4638,a4640,a4642,a4644,a4646,a4648,a4650,
a4652,a4654,a4656,a4658,a4660,a4662,a4664,a4666,a4668,a4670,a4672,a4674,a4676,a4678,a4680,
a4682,a4684,a4686,a4688,a4690,a4692,a4694,a4696,a4698,a4700,a4702,a4704,a4706,a4708,a4710,
a4712,a4714,a4716,a4718,a4720,a4722,a4724,a4726,a4728,a4730,a4732,a4734,a4736,a4738,a4740,
a4742,a4744,a4746,a4748,a4750,a4752,a4754,a4756,a4758,a4760,a4762,a4764,a4766,a4768,a4770,
a4772,a4774,a4776,a4778,a4780,a4782,a4784,a4786,a4788,a4790,a4792,a4794,a4796,a4798,a4800,
a4802,a4804,a4806,a4808,a4810,a4812,a4814,a4816,a4818,a4820,a4822,a4824,a4826,a4828,a4830,
a4832,a4834,a4836,a4838,a4840,a4842,a4844,a4846,a4848,a4850,a4852,a4854,a4856,a4858,a4860,
a4862,a4864,a4866,a4868,a4870,a4872,a4874,a4876,a4878,a4880,a4882,a4884,a4886,a4888,a4890,
a4892,a4894,a4896,a4898,a4900,a4902,a4904,a4906,a4908,a4910,a4912,a4914,a4916,a4918,a4920,
a4922,a4924,a4926,a4928,a4930,a4932,a4934,a4936,a4938,a4940,a4942,a4944,a4946,a4948,a4950,
a4952,a4954,a4956,a4958,a4960,a4962,a4964,a4966,a4968,a4970,a4972,a4974,a4976,a4978,a4980,
a4982,a4984,a4986,a4988,a4990,a4992,a4994,a4996,a4998,a5000,a5002,a5004,a5006,a5008,a5010,
a5012,a5014,a5016,a5018,a5020,a5022,a5024,a5026,a5028,a5030,a5032,a5034,a5036,a5038,a5040,
a5042,a5044,a5046,a5048,a5050,a5052,a5054,a5056,a5058,a5060,a5062,a5064,a5066,a5068,a5070,
a5072,a5074,a5076,a5078,a5080,a5082,a5084,a5086,a5088,a5090,a5092,a5094,a5096,a5098,a5100,
a5102,a5104,a5106,a5108,a5110,a5112,a5114,a5116,a5118,a5120,a5122,a5124,a5126,a5128,a5130,
a5132,a5134,a5136,a5138,a5140,a5142,a5144,a5146,a5148,a5150,a5152,a5154,a5156,a5158,a5160,
a5162,a5164,a5166,a5168,a5170,a5172,a5174,a5176,a5178,a5180,a5182,a5184,a5186,a5188,a5190,
a5192,a5194,a5196,a5198,a5200,a5202,a5204,a5206,a5208,a5210,a5212,a5214,a5216,a5218,a5220,
a5222,a5224,a5226,a5228,a5230,a5232,a5234,a5236,a5238,a5240,a5242,a5244,a5246,a5248,a5250,
a5252,a5254,a5256,a5258,a5260,a5262,a5264,a5266,a5268,a5270,a5272,a5274,a5276,a5278,a5280,
a5282,a5284,a5286,a5288,a5290,a5292,a5294,a5296,a5298,a5300,a5302,a5304,a5306,a5308,a5310,
a5312,a5314,a5316,a5318,a5320,a5322,a5324,a5326,a5328,a5330,a5332,a5334,a5336,a5338,a5340,
a5342,a5344,a5346,a5348,a5350,a5352,a5354,a5356,a5358,a5360,a5362,a5364,a5366,a5368,a5370,
a5372,a5374,a5376,a5378,a5380,a5382,a5384,a5386,a5388,a5390,a5392,a5394,a5396,a5398,a5400,
a5402,a5404,a5406,a5408,a5410,a5412,a5414,a5416,a5418,a5420,a5422,a5424,a5426,a5428,a5430,
a5432,a5434,a5436,a5438,a5440,a5442,a5444,a5446,a5448,a5450,a5452,a5454,a5456,a5458,a5460,
a5462,a5464,a5466,a5468,a5470,a5472,a5474,a5476,a5478,a5480,a5482,a5484,a5486,a5488,a5490,
a5492,a5494,a5496,a5498,a5500,a5502,a5504,a5506,a5508,a5510,a5512,a5514,a5516,a5518,a5520,
a5522,a5524,a5526,a5528,a5530,a5532,a5534,a5536,a5538,a5540,a5542,a5544,a5546,a5548,a5550,
a5552,a5554,a5556,a5558,a5560,a5562,a5564,a5566,a5568,a5570,a5572,a5574,a5576,a5578,a5580,
a5582,a5584,a5586,a5588,a5590,a5592,a5594,a5596,a5598,a5600,a5602,a5604,a5606,a5608,a5610,
a5612,a5614,a5616,a5618,a5620,a5622,a5624,a5626,a5628,a5630,a5632,a5634,a5636,a5638,a5640,
a5642,a5644,a5646,a5648,a5650,a5652,a5654,a5656,a5658,a5660,a5662,a5664,a5666,a5668,a5670,
a5672,a5674,a5676,a5678,a5680,a5682,a5684,a5686,a5688,a5690,a5692,a5694,a5696,a5698,a5700,
a5702,a5704,a5706,a5708,a5710,a5712,a5714,a5716,a5718,a5720,a5722,a5724,a5726,a5728,a5730,
a5732,a5734,a5736,a5738,a5740,a5742,a5744,a5746,a5748,a5750,a5752,a5754,a5756,a5758,a5760,
a5762,a5764,a5766,a5768,a5770,a5772,a5774,a5776,a5778,a5780,a5782,a5784,a5786,a5788,a5790,
a5792,a5794,a5796,a5798,a5800,a5802,a5804,a5806,a5808,a5810,a5812,a5814,a5816,a5818,a5820,
a5822,a5824,a5826,a5828,a5830,a5832,a5834,a5836,a5838,a5840,a5842,a5844,a5846,a5848,a5850,
a5852,a5854,a5856,a5858,a5860,a5862,a5864,a5866,a5868,a5870,a5872,a5874,a5876,a5878,a5880,
a5882,a5884,a5886,a5888,a5890,a5892,a5894,a5896,a5898,a5900,a5902,a5904,a5906,a5908,a5910,
a5912,a5914,a5916,a5918,a5920,a5922,a5924,a5926,a5928,a5930,a5932,a5934,a5936,a5938,a5940,
a5942,a5944,a5946,a5948,a5950,a5952,a5954,a5956,a5958,a5960,a5962,a5964,a5966,a5968,a5970,
a5972,a5974,a5976,a5978,a5980,a5982,a5984,a5986,a5988,a5990,a5992,a5994,a5996,a5998,a6000,
a6002,a6004,a6006,a6008,a6010,a6012,a6014,a6016,a6018,a6020,a6022,a6024,a6026,a6028,a6030,
a6032,a6034,a6036,a6038,a6040,a6042,a6044,a6046,a6048,a6050,a6052,a6054,a6056,a6058,a6060,
a6062,a6064,a6066,a6068,a6070,a6072,a6074,a6076,a6078,a6080,a6082,a6084,a6086,a6088,a6090,
a6092,a6094,a6096,a6098,a6100,a6102,a6104,a6106,a6108,a6110,a6112,a6114,a6116,a6118,a6120,
a6122,a6124,a6126,a6128,a6130,a6132,a6134,a6136,a6138,a6140,a6142,a6144,a6146,a6148,a6150,
a6152,a6154,a6156,a6158,a6160,a6162,a6164,a6166,a6168,a6170,a6172,a6174,a6176,a6178,a6180,
a6182,a6184,a6186,a6188,a6190,a6192,a6194,a6196,a6198,a6200,a6202,a6204,a6206,a6208,a6210,
a6212,a6214,a6216,a6218,a6220,a6222,a6224,a6226,a6228,a6230,a6232,a6234,a6236,a6238,a6240,
a6242,a6244,a6246,a6248,a6250,a6252,a6254,a6256,a6258,a6260,a6262,a6264,a6266,a6268,a6270,
a6272,a6274,a6276,a6278,a6280,a6282,a6284,a6286,a6288,a6290,a6292,a6294,a6296,a6298,a6300,
a6302,a6304,a6306,a6308,a6310,a6312,a6314,a6316,a6318,a6320,a6322,a6324,a6326,a6328,a6330,
a6332,a6334,a6336,a6338,a6340,a6342,a6344,a6346,a6348,a6350,a6352,a6354,a6356,a6358,a6360,
a6362,a6364,a6366,a6368,a6370,a6372,a6374,a6376,a6378,a6380,a6382,a6384,a6386,a6388,a6390,
a6392,a6394,a6396,a6398,a6400,a6402,a6404,a6406,a6408,a6410,a6412,a6414,a6416,a6418,a6420,
a6422,a6424,a6426,a6428,a6430,a6432,a6434,a6436,a6438,a6440,a6442,a6444,a6446,a6448,a6450,
a6452,a6454,a6456,a6458,a6460,a6462,a6464,a6466,a6468,a6470,a6472,a6474,a6476,a6478,a6480,
a6482,a6484,a6486,a6488,a6490,a6492,a6494,a6496,a6498,a6500,a6502,a6504,a6506,a6508,a6510,
a6512,a6514,a6516,a6518,a6520,a6522,a6524,a6526,a6528,a6530,a6532,a6534,a6536,a6538,a6540,
a6542,a6544,a6546,a6548,a6550,a6552,a6554,a6556,a6558,a6560,a6562,a6564,a6566,a6568,a6570,
a6572,a6574,a6576,a6578,a6580,a6582,a6584,a6586,a6588,a6590,a6592,a6594,a6596,a6598,a6600,
a6602,a6604,a6606,a6608,a6610,a6612,a6614,a6616,a6618,a6620,a6622,a6624,a6626,a6628,a6630,
a6632,a6634,a6636,a6638,a6640,a6642,a6644,a6646,a6648,a6650,a6652,a6654,a6656,a6658,a6660,
a6662,a6664,a6666,a6668,a6670,a6672,a6674,a6676,a6678,a6680,a6682,a6684,a6686,a6688,a6690,
a6692,a6694,a6696,a6698,a6700,a6702,a6704,a6706,a6708,a6710,a6712,a6714,a6716,a6718,a6720,
a6722,a6724,a6726,a6728,a6730,a6732,a6734,a6736,a6738,a6740,a6742,a6744,a6746,a6748,a6750,
a6752,a6754,a6756,a6758,a6760,a6762,a6764,a6766,a6768,a6770,a6772,a6774,a6776,a6778,a6780,
a6782,a6784,a6786,a6788,a6790,a6792,a6794,a6796,a6798,a6800,a6802,a6804,a6806,a6808,a6810,
a6812,a6814,a6816,a6818,a6820,a6822,a6824,a6826,a6828,a6830,a6832,a6834,a6836,a6838,a6840,
a6842,a6844,a6846,a6848,a6850,a6852,a6854,a6856,a6858,a6860,a6862,a6864,a6866,a6868,a6870,
a6872,a6874,a6876,a6878,a6880,a6882,a6884,a6886,a6888,a6890,a6892,a6894,a6896,a6898,a6900,
a6902,a6904,a6906,a6908,a6910,a6912,a6914,a6916,a6918,a6920,a6922,a6924,a6926,a6928,a6930,
a6932,a6934,a6936,a6938,a6940,a6942,a6944,a6946,a6948,a6950,a6952,a6954,a6956,a6958,a6960,
a6962,a6964,a6966,a6968,a6970,a6972,a6974,a6976,a6978,a6980,a6982,a6984,a6986,a6988,a6990,
a6992,a6994,a6996,a6998,a7000,a7002,a7004,a7006,a7008,a7010,a7012,a7014,a7016,a7018,a7020,
a7022,a7024,a7026,a7028,a7030,a7032,a7034,a7036,a7038,a7040,a7042,a7044,a7046,a7048,a7050,
a7052,a7054,a7056,a7058,a7060,a7062,a7064,a7066,a7068,a7070,a7072,a7074,a7076,a7078,a7080,
a7082,a7084,a7086,a7088,a7090,a7092,a7094,a7096,a7098,a7100,a7102,a7104,a7106,a7108,a7110,
a7112,a7114,a7116,a7118,a7120,a7122,a7124,a7126,a7128,a7130,a7132,a7134,a7136,a7138,a7140,
a7142,a7144,a7146,a7148,a7150,a7152,a7154,a7156,a7158,a7160,a7162,a7164,a7166,a7168,a7170,
a7172,a7174,a7176,a7178,a7180,a7182,a7184,a7186,a7188,a7190,a7192,a7194,a7196,a7198,a7200,
a7202,a7204,a7206,a7208,a7210,a7212,a7214,a7216,a7218,a7220,a7222,a7224,a7226,a7228,a7230,
a7232,a7234,a7236,a7238,a7240,a7242,a7244,a7246,a7248,a7250,a7252,a7254,a7256,a7258,a7260,
a7262,a7264,a7266,a7268,a7270,a7272,a7274,a7276,a7278,a7280,a7282,a7284,a7286,a7288,a7290,
a7292,a7294,a7296,a7298,a7300,a7302,a7304,a7306,a7308,a7310,a7312,a7314,a7316,a7318,a7320,
a7322,a7324,a7326,a7328,a7330,a7332,a7334,a7336,a7338,a7340,a7342,a7344,a7346,a7348,a7350,
a7352,a7354,a7356,a7358,a7360,a7362,a7364,a7366,a7368,a7370,a7372,a7374,a7376,a7378,a7380,
a7382,a7384,a7386,a7388,a7390,a7392,a7394,a7396,a7398,a7400,a7402,a7404,a7406,a7408,a7410,
a7412,a7414,a7416,a7418,a7420,a7422,a7424,a7426,a7428,a7430,a7432,a7434,a7436,a7438,a7440,
a7442,a7444,a7446,a7448,a7450,a7452,a7454,a7456,a7458,a7460,a7462,a7464,a7466,a7468,a7470,
a7472,a7474,a7476,a7478,a7480,a7482,a7484,a7486,a7488,a7490,a7492,a7494,a7496,a7498,a7500,
a7502,a7504,a7506,a7508,a7510,a7512,a7514,a7516,a7518,a7520,a7522,a7524,a7526,a7528,a7530,
a7532,a7534,a7536,a7538,a7540,a7542,a7544,a7546,a7548,a7550,a7552,a7554,a7556,a7558,a7560,
a7562,a7564,a7566,a7568,a7570,a7572,a7574,a7576,a7578,a7580,a7582,a7584,a7586,a7588,a7590,
a7592,a7594,a7596,a7598,a7600,a7602,a7604,a7606,a7608,a7610,a7612,a7614,a7616,a7618,a7620,
a7622,a7624,a7626,a7628,a7630,a7632,a7634,a7636,a7638,a7640,a7642,a7644,a7646,a7648,a7650,
a7652,a7654,a7656,a7658,a7660,a7662,a7664,a7666,a7668,a7670,a7672,a7674,a7676,a7678,a7680,
a7682,a7684,a7686,a7688,a7690,a7692,a7694,a7696,a7698,a7700,a7702,a7704,a7706,a7708,a7710,
a7712,a7714,a7716,a7718,a7720,a7722,a7724,a7726,a7728,a7730,a7732,a7734,a7736,a7738,a7740,
a7742,a7744,a7746,a7748,a7750,a7752,a7754,a7756,a7758,a7760,a7762,a7764,a7766,a7768,a7770,
a7772,a7774,a7776,a7778,a7780,a7782,a7784,a7786,a7788,a7790,a7792,a7794,a7796,a7798,a7800,
a7802,a7804,a7806,a7808,a7810,a7812,a7814,a7816,a7818,a7820,a7822,a7824,a7826,a7828,a7830,
a7832,a7834,a7836,a7838,a7840,a7842,a7844,a7846,a7848,a7850,a7852,a7854,a7856,a7858,a7860,
a7862,a7864,a7866,a7868,a7870,a7872,a7874,a7876,a7878,a7880,a7882,a7884,a7886,a7888,a7890,
a7892,a7894,a7896,a7898,a7900,a7902,a7904,a7906,a7908,a7910,a7912,a7914,a7916,a7918,a7920,
a7922,a7924,a7926,a7928,a7930,a7932,a7934,a7936,a7938,a7940,a7942,a7944,a7946,a7948,a7950,
a7952,a7954,a7956,a7958,a7960,a7962,a7964,a7966,a7968,a7970,a7972,a7974,a7976,a7978,a7980,
a7982,a7984,a7986,a7988,a7990,a7992,a7994,a7996,a7998,a8000,a8002,a8004,a8006,a8008,a8010,
a8012,a8014,a8016,a8018,a8020,a8022,a8024,a8026,a8028,a8030,a8032,a8034,a8036,a8038,a8040,
a8042,a8044,a8046,a8048,a8050,a8052,a8054,a8056,a8058,a8060,a8062,a8064,a8066,a8068,a8070,
a8072,a8074,a8076,a8078,a8080,a8082,a8084,a8086,a8088,a8090,a8092,a8094,a8096,a8098,a8100,
a8102,a8104,a8106,a8108,a8110,a8112,a8114,a8116,a8118,a8120,a8122,a8124,a8126,a8128,a8130,
a8132,a8134,a8136,a8138,a8140,a8142,a8144,a8146,a8148,a8150,a8152,a8154,a8156,a8158,a8160,
a8162,a8164,a8166,a8168,a8170,a8172,a8174,a8176,a8178,a8180,a8182,a8184,a8186,a8188,a8190,
a8192,a8194,a8196,a8198,a8200,a8202,a8204,a8206,a8208,a8210,a8212,a8214,a8216,a8218,a8220,
a8222,a8224,a8226,a8228,a8230,a8232,a8234,a8236,a8238,a8240,a8242,a8244,a8246,a8248,a8250,
a8252,a8254,a8256,a8258,a8260,a8262,a8264,a8266,a8268,a8270,a8272,a8274,a8276,a8278,a8280,
a8282,a8284,a8286,a8288,a8290,a8292,a8294,a8296,a8298,a8300,a8302,a8304,a8306,a8308,a8310,
a8312,a8314,a8316,a8318,a8320,a8322,a8324,a8326,a8328,a8330,a8332,a8334,a8336,a8338,a8340,
a8342,a8344,a8346,a8348,a8350,a8352,a8354,a8356,a8358,a8360,a8362,a8364,a8366,a8368,a8370,
a8372,a8374,a8376,a8378,a8380,a8382,a8384,a8386,a8388,a8390,a8392,a8394,a8396,a8398,a8400,
a8402,a8404,a8406,a8408,a8410,a8412,a8414,a8416,a8418,a8420,a8422,a8424,a8426,a8428,a8430,
a8432,a8434,a8436,a8438,a8440,a8442,a8444,a8446,a8448,a8450,a8452,a8454,a8456,a8458,a8460,
a8462,a8464,a8466,a8468,a8470,a8472,a8474,a8476,a8478,a8480,a8482,a8484,a8486,a8488,a8490,
a8492,a8494,a8496,a8498,a8500,a8502,a8504,a8506,a8508,a8510,a8512,a8514,a8516,a8518,a8520,
a8522,a8524,a8526,a8528,a8530,a8532,a8534,a8536,a8538,a8540,a8542,a8544,a8546,a8548,a8550,
a8552,a8554,a8556,a8558,a8560,a8562,a8564,a8566,a8568,a8570,a8572,a8574,a8576,a8578,a8580,
a8582,a8584,a8586,a8588,a8590,a8592,a8594,a8596,a8598,a8600,a8602,a8604,a8606,a8608,a8610,
a8612,a8614,a8616,a8618,a8620,a8622,a8624,a8626,a8628,a8630,a8632,a8634,a8636,a8638,a8640,
a8642,a8644,a8646,a8648,a8650,a8652,a8654,a8656,a8658,a8660,a8662,a8664,a8666,a8668,a8670,
a8672,a8674,a8676,a8678,a8680,a8682,a8684,a8686,a8688,a8690,a8692,a8694,a8696,a8698,a8700,
a8702,a8704,a8706,a8708,a8710,a8712,a8714,a8716,a8718,a8720,a8722,a8724,a8726,a8728,a8730,
a8732,a8734,a8736,a8738,a8740,a8742,a8744,a8746,a8748,a8750,a8752,a8754,a8756,a8758,a8760,
a8762,a8764,a8766,a8768,a8770,a8772,a8774,a8776,a8778,a8780,a8782,a8784,a8786,a8788,a8790,
a8792,a8794,a8796,a8798,a8800,a8802,a8804,a8806,a8808,a8810,a8812,a8814,a8816,a8818,a8820,
a8822,a8824,a8826,a8828,a8830,a8832,a8834,a8836,a8838,a8840,a8842,a8844,a8846,a8848,a8850,
a8852,a8854,a8856,a8858,a8860,a8862,a8864,a8866,a8868,a8870,a8872,a8874,a8876,a8878,a8880,
a8882,a8884,a8886,a8888,a8890,a8892,a8894,a8896,a8898,a8900,a8902,a8904,a8906,a8908,a8910,
a8912,a8914,a8916,a8918,a8920,a8922,a8924,a8926,a8928,a8930,a8932,a8934,a8936,a8938,a8940,
a8942,a8944,a8946,a8948,a8950,a8952,a8954,a8956,a8958,a8960,a8962,a8964,a8966,a8968,a8970,
a8972,a8974,a8976,a8978,a8980,a8982,a8984,a8986,a8988,a8990,a8992,a8994,a8996,a8998,a9000,
a9002,a9004,a9006,a9008,a9010,a9012,a9014,a9016,a9018,a9020,a9022,a9024,a9026,a9028,a9030,
a9032,a9034,a9036,a9038,a9040,a9042,a9044,a9046,a9048,a9050,a9052,a9054,a9056,a9058,a9060,
a9062,a9064,a9066,a9068,a9070,a9072,a9074,a9076,a9078,a9080,a9082,a9084,a9086,a9088,a9090,
a9092,a9094,a9096,a9098,a9100,a9102,a9104,a9106,a9108,a9110,a9112,a9114,a9116,a9118,a9120,
a9122,a9124,a9126,a9128,a9130,a9132,a9134,a9136,a9138,a9140,a9142,a9144,a9146,a9148,a9150,
a9152,a9154,a9156,a9158,a9160,a9162,a9164,a9166,a9168,a9170,a9172,a9174,a9176,a9178,a9180,
a9182,a9184,a9186,a9188,a9190,a9192,a9194,a9196,a9198,a9200,a9202,a9204,a9206,a9208,a9210,
a9212,a9214,a9216,a9218,a9220,a9222,a9224,a9226,a9228,a9230,a9232,a9234,a9236,a9238,a9240,
a9242,a9244,a9246,a9248,a9250,a9252,a9254,a9256,a9258,a9260,a9262,a9264,a9266,a9268,a9270,
a9272,a9274,a9276,a9278,a9280,a9282,a9284,a9286,a9288,a9290,a9292,a9294,a9296,a9298,a9300,
a9302,a9304,a9306,a9308,a9310,a9312,a9314,a9316,a9318,a9320,a9322,a9324,a9326,a9328,a9330,
a9332,a9334,a9336,a9338,a9340,a9342,a9344,a9346,a9348,a9350,a9352,a9354,a9356,a9358,a9360,
a9362,a9364,a9366,a9368,a9370,a9372,a9374,a9376,a9378,a9380,a9382,a9384,a9386,a9388,a9390,
a9392,a9394,a9396,a9398,a9400,a9402,a9404,a9406,a9408,a9410,a9412,a9414,a9416,a9418,a9420,
a9422,a9424,a9426,a9428,a9430,a9432,a9434,a9436,a9438,a9440,a9442,a9444,a9446,a9448,a9450,
a9452,a9454,a9456,a9458,a9460,a9462,a9464,a9466,a9468,a9470,a9472,a9474,a9476,a9478,a9480,
a9482,a9484,a9486,a9488,a9490,a9492,a9494,a9496,a9498,a9500,a9502,a9504,a9506,a9508,a9510,
a9512,a9514,a9516,a9518,a9520,a9522,a9524,a9526,a9528,a9530,a9532,a9534,a9536,a9538,a9540,
a9542,a9544,a9546,a9548,a9550,a9552,a9554,a9556,a9558,a9560,a9562,a9564,a9566,a9568,a9570,
a9572,a9574,a9576,a9578,a9580,a9582,a9584,a9586,a9588,a9590,a9592,a9594,a9596,a9598,a9600,
a9602,a9604,a9606,a9608,a9610,a9612,a9614,a9616,a9618,a9620,a9622,a9624,a9626,a9628,a9630,
a9632,a9634,a9636,a9638,a9640,a9642,a9644,a9646,a9648,a9650,a9652,a9654,a9656,a9658,a9660,
a9662,a9664,a9666,a9668,a9670,a9672,a9674,a9676,a9678,a9680,a9682,a9684,a9686,a9688,a9690,
a9692,a9694,a9696,a9698,a9700,a9702,a9704,a9706,a9708,a9710,a9712,a9714,a9716,a9718,a9720,
a9722,a9724,a9726,a9728,a9730,a9732,a9734,a9736,a9738,a9740,a9742,a9744,a9746,a9748,a9750,
a9752,a9754,a9756,a9758,a9760,a9762,a9764,a9766,a9768,a9770,a9772,a9774,a9776,a9778,a9780,
a9782,a9784,a9786,a9788,a9790,a9792,a9794,a9796,a9798,a9800,a9802,a9804,a9806,a9808,a9810,
a9812,a9814,a9816,a9818,a9820,a9822,a9824,a9826,a9828,a9830,a9832,a9834,a9836,a9838,a9840,
a9842,a9844,a9846,a9848,a9850,a9852,a9854,a9856,a9858,a9860,a9862,a9864,a9866,a9868,a9870,
a9872,a9874,a9876,a9878,a9880,a9882,a9884,a9886,a9888,a9890,a9892,a9894,a9896,a9898,a9900,
a9902,a9904,a9906,a9908,a9910,a9912,a9914,a9916,a9918,a9920,a9922,a9924,a9926,a9928,a9930,
a9932,a9934,a9936,a9938,a9940,a9942,a9944,a9946,a9948,a9950,a9952,a9954,a9956,a9958,a9960,
a9962,a9964,a9966,a9968,a9970,a9972,a9974,a9976,a9978,a9980,a9982,a9984,a9986,a9988,a9990,
a9992,a9994,a9996,a9998,a10000,a10002,a10004,a10006,a10008,a10010,a10012,a10014,a10016,a10018,a10020,
a10022,a10024,a10026,a10028,a10030,a10032,a10034,a10036,a10038,a10040,a10042,a10044,a10046,a10048,a10050,
a10052,a10054,a10056,a10058,a10060,a10062,a10064,a10066,a10068,a10070,a10072,a10074,a10076,a10078,a10080,
a10082,a10084,a10086,a10088,a10090,a10092,a10094,a10096,a10098,a10100,a10102,a10104,a10106,a10108,a10110,
a10112,a10114,a10116,a10118,a10120,a10122,a10124,a10126,a10128,a10130,a10132,a10134,a10136,a10138,a10140,
a10142,a10144,a10146,a10148,a10150,a10152,a10154,a10156,a10158,a10160,a10162,a10164,a10166,a10168,a10170,
a10172,a10174,a10176,a10178,a10180,a10182,a10184,a10186,a10188,a10190,a10192,a10194,a10196,a10198,a10200,
a10202,a10204,a10206,a10208,a10210,a10212,a10214,a10216,a10218,a10220,a10222,a10224,a10226,a10228,a10230,
a10232,a10234,a10236,a10238,a10240,a10242,a10244,a10246,a10248,a10250,a10252,a10254,a10256,a10258,a10260,
a10262,a10264,a10266,a10268,a10270,a10272,a10274,a10276,a10278,a10280,a10282,a10284,a10286,a10288,a10290,
a10292,a10294,a10296,a10298,a10300,a10302,a10304,a10306,a10308,a10310,a10312,a10314,a10316,a10318,a10320,
a10322,a10324,a10326,a10328,a10330,a10332,a10334,a10336,a10338,a10340,a10342,a10344,a10346,a10348,a10350,
a10352,a10354,a10356,a10358,a10360,a10362,a10364,a10366,a10368,a10370,a10372,a10374,a10376,a10378,a10380,
a10382,a10384,a10386,a10388,a10390,a10392,a10394,a10396,a10398,a10400,a10402,a10404,a10406,a10408,a10410,
a10412,a10414,a10416,a10418,a10420,a10422,a10424,a10426,a10428,a10430,a10432,a10434,a10436,a10438,a10440,
a10442,a10444,a10446,a10448,a10450,a10452,a10454,a10456,a10458,a10460,a10462,a10464,a10466,a10468,a10470,
a10472,a10474,a10476,a10478,a10480,a10482,a10484,a10486,a10488,a10490,a10492,a10494,a10496,a10498,a10500,
a10502,a10504,a10506,a10508,a10510,a10512,a10514,a10516,a10518,a10520,a10522,a10524,a10526,a10528,a10530,
a10532,a10534,a10536,a10538,a10540,a10542,a10544,a10546,a10548,a10550,a10552,a10554,a10556,a10558,a10560,
a10562,a10564,a10566,a10568,a10570,a10572,a10574,a10576,a10578,a10580,a10582,a10584,a10586,a10588,a10590,
a10592,a10594,a10596,a10598,a10600,a10602,a10604,a10606,a10608,a10610,a10612,a10614,a10616,a10618,a10620,
a10622,a10624,a10626,a10628,a10630,a10632,a10634,a10636,a10638,a10640,a10642,a10644,a10646,a10648,a10650,
a10652,a10654,a10656,a10658,a10660,a10662,a10664,a10666,a10668,a10670,a10672,a10674,a10676,a10678,a10680,
a10682,a10684,a10686,a10688,a10690,a10692,a10694,a10696,a10698,a10700,a10702,a10704,a10706,a10708,a10710,
a10712,a10714,a10716,a10718,a10720,a10722,a10724,a10726,a10728,a10730,a10732,a10734,a10736,a10738,a10740,
a10742,a10744,a10746,a10748,a10750,a10752,a10754,a10756,a10758,a10760,a10762,a10764,a10766,a10768,a10770,
a10772,a10774,a10776,a10778,a10780,a10782,a10784,a10786,a10788,a10790,a10792,a10794,a10796,a10798,a10800,
a10802,a10804,a10806,a10808,a10810,a10812,a10814,a10816,a10818,a10820,a10822,a10824,a10826,a10828,a10830,
a10832,a10834,a10836,a10838,a10840,a10842,a10844,a10846,a10848,a10850,a10852,a10854,a10856,a10858,a10860,
a10862,a10864,a10866,a10868,a10870,a10872,a10874,a10876,a10878,a10880,a10882,a10884,a10886,a10888,a10890,
a10892,a10894,a10896,a10898,a10900,a10902,a10904,a10906,a10908,a10910,a10912,a10914,a10916,a10918,a10920,
a10922,a10924,a10926,a10928,a10930,a10932,a10934,a10936,a10938,a10940,a10942,a10944,a10946,a10948,a10950,
a10952,a10954,a10956,a10958,a10960,a10962,a10964,a10966,a10968,a10970,a10972,a10974,a10976,a10978,a10980,
a10982,a10984,a10986,a10988,a10990,a10992,a10994,a10996,a10998,a11000,a11002,a11004,a11006,a11008,a11010,
a11012,a11014,a11016,a11018,a11020,a11022,a11024,a11026,a11028,a11030,a11032,a11034,a11036,a11038,a11040,
a11042,a11044,a11046,a11048,a11050,a11052,a11054,a11056,a11058,a11060,a11062,a11064,a11066,a11068,a11070,
a11072,a11074,a11076,a11078,a11080,a11082,a11084,a11086,a11088,a11090,a11092,a11094,a11096,a11098,a11100,
a11102,a11104,a11106,a11108,a11110,a11112,a11114,a11116,a11118,a11120,a11122,a11124,a11126,a11128,a11130,
a11132,a11134,a11136,a11138,a11140,a11142,a11144,a11146,a11148,a11150,a11152,a11154,a11156,a11158,a11160,
a11162,a11164,a11166,a11168,a11170,a11172,a11174,a11176,a11178,a11180,a11182,a11184,a11186,a11188,a11190,
a11192,a11194,a11196,a11198,a11200,a11202,a11204,a11206,a11208,a11210,a11212,a11214,a11216,a11218,a11220,
a11222,a11224,a11226,a11228,a11230,a11232,a11234,a11236,a11238,a11240,a11242,a11244,a11246,a11248,a11250,
a11252,a11254,a11256,a11258,a11260,a11262,a11264,a11266,a11268,a11270,a11272,a11274,a11276,a11278,a11280,
a11282,a11284,a11286,a11288,a11290,a11292,a11294,a11296,a11298,a11300,a11302,a11304,a11306,a11308,a11310,
a11312,a11314,a11316,a11318,a11320,a11322,a11324,a11326,a11328,a11330,a11332,a11334,a11336,a11338,a11340,
a11342,a11344,a11346,a11348,a11350,a11352,a11354,a11356,a11358,a11360,a11362,a11364,a11366,a11368,a11370,
a11372,a11374,a11376,a11378,a11380,a11382,a11384,a11386,a11388,a11390,a11392,a11394,a11396,a11398,a11400,
a11402,a11404,a11406,a11408,a11410,a11412,a11414,a11416,a11418,a11420,a11422,a11424,a11426,a11428,a11430,
a11432,a11434,a11436,a11438,a11440,a11442,a11444,a11446,a11448,a11450,a11452,a11454,a11456,a11458,a11460,
a11462,a11464,a11466,a11468,a11470,a11472,a11474,a11476,a11478,a11480,a11482,a11484,a11486,a11488,a11490,
a11492,a11494,a11496,a11498,a11500,a11502,a11504,a11506,a11508,a11510,a11512,a11514,a11516,a11518,a11520,
a11522,a11524,a11526,a11528,a11530,a11532,a11534,a11536,a11538,a11540,a11542,a11544,a11546,a11548,a11550,
a11552,a11554,a11556,a11558,a11560,a11562,a11564,a11566,a11568,a11570,a11572,a11574,a11576,a11578,a11580,
a11582,a11584,a11586,a11588,a11590,a11592,a11594,a11596,a11598,a11600,a11602,a11604,a11606,a11608,a11610,
a11612,a11614,a11616,a11618,a11620,a11622,a11624,a11626,a11628,a11630,a11632,a11634,a11636,a11638,a11640,
a11642,a11644,a11646,a11648,a11650,a11652,a11654,a11656,a11658,a11660,a11662,a11664,a11666,a11668,a11670,
a11672,a11674,a11676,a11678,a11680,a11682,a11684,a11686,a11688,a11690,a11692,a11694,a11696,a11698,a11700,
a11702,a11704,a11706,a11708,a11710,a11712,a11714,a11716,a11718,a11720,a11722,a11724,a11726,a11728,a11730,
a11732,a11734,a11736,a11738,a11740,a11742,a11744,a11746,a11748,a11750,a11752,a11754,a11756,a11758,a11760,
a11762,a11764,a11766,a11768,a11770,a11772,a11774,a11776,a11778,a11780,a11782,a11784,a11786,a11788,a11790,
a11792,a11794,a11796,a11798,a11800,a11802,a11804,a11806,a11808,a11810,a11812,a11814,a11816,a11818,a11820,
a11822,a11824,a11826,a11828,a11830,a11832,a11834,a11836,a11838,a11840,a11842,a11844,a11846,a11848,a11850,
a11852,a11854,a11856,a11858,a11860,a11862,a11864,a11866,a11868,a11870,a11872,a11874,a11876,a11878,a11880,
a11882,a11884,a11886,a11888,a11890,a11892,a11894,a11896,a11898,a11900,a11902,a11904,a11906,a11908,a11910,
a11912,a11914,a11916,a11918,a11920,a11922,a11924,a11926,a11928,a11930,a11932,a11934,a11936,a11938,a11940,
a11942,a11944,a11946,a11948,a11950,a11952,a11954,a11956,a11958,a11960,a11962,a11964,a11966,a11968,a11970,
a11972,a11974,a11976,a11978,a11980,a11982,a11984,a11986,a11988,a11990,a11992,a11994,a11996,a11998,a12000,
a12002,a12004,a12006,a12008,a12010,a12012,a12014,a12016,a12018,a12020,a12022,a12024,a12026,a12028,a12030,
a12032,a12034,a12036,a12038,a12040,a12042,a12044,a12046,a12048,a12050,a12052,a12054,a12056,a12058,a12060,
a12062,a12064,a12066,a12068,a12070,a12072,a12074,a12076,a12078,a12080,a12082,a12084,a12086,a12088,a12090,
a12092,a12094,a12096,a12098,a12100,a12102,a12104,a12106,a12108,a12110,a12112,a12114,a12116,a12118,a12120,
a12122,a12124,a12126,a12128,a12130,a12132,a12134,a12136,a12138,a12140,a12142,a12144,a12146,a12148,a12150,
a12152,a12154,a12156,a12158,a12160,a12162,a12164,a12166,a12168,a12170,a12172,a12174,a12176,a12178,a12180,
a12182,a12184,a12186,a12188,a12190,a12192,a12194,a12196,a12198,a12200,a12202,a12204,a12206,a12208,a12210,
a12212,a12214,a12216,a12218,a12220,a12222,a12224,a12226,a12228,a12230,a12232,a12234,a12236,a12238,a12240,
a12242,a12244,a12246,a12248,a12250,a12252,a12254,a12256,a12258,a12260,a12262,a12264,a12266,a12268,a12270,
a12272,a12274,a12276,a12278,a12280,a12282,a12284,a12286,a12288,a12290,a12292,a12294,a12296,a12298,a12300,
a12302,a12304,a12306,a12308,a12310,a12312,a12314,a12316,a12318,a12320,a12322,a12324,a12326,a12328,a12330,
a12332,a12334,a12336,a12338,a12340,a12342,a12344,a12346,a12348,a12350,a12352,a12354,a12356,a12358,a12360,
a12362,a12364,a12366,a12368,a12370,a12372,a12374,a12376,a12378,a12380,a12382,a12384,a12386,a12388,a12390,
a12392,a12394,a12396,a12398,a12400,a12402,a12404,a12406,a12408,a12410,a12412,a12414,a12416,a12418,a12420,
a12422,a12424,a12426,a12428,a12430,a12432,a12434,a12436,a12438,a12440,a12442,a12444,a12446,a12448,a12450,
a12452,a12454,a12456,a12458,a12460,a12462,a12464,a12466,a12468,a12470,a12472,a12474,a12476,a12478,a12480,
a12482,a12484,a12486,a12488,a12490,a12492,a12494,a12496,a12498,a12500,a12502,a12504,a12506,a12508,a12510,
a12512,a12514,a12516,a12518,a12520,a12522,a12524,a12526,a12528,a12530,a12532,a12534,a12536,a12538,a12540,
a12542,a12544,a12546,a12548,a12550,a12552,a12554,a12556,a12558,a12560,a12562,a12564,a12566,a12568,a12570,
a12572,a12574,a12576,a12578,a12580,a12582,a12584,a12586,a12588,a12590,a12592,a12594,a12596,a12598,a12600,
a12602,a12604,a12606,a12608,a12610,a12612,a12614,a12616,a12618,a12620,a12622,a12624,a12626,a12628,a12630,
a12632,a12634,a12636,a12638,a12640,a12642,a12644,a12646,a12648,a12650,a12652,a12654,a12656,a12658,a12660,
a12662,a12664,a12666,a12668,a12670,a12672,a12674,a12676,a12678,a12680,a12682,a12684,a12686,a12688,a12690,
a12692,a12694,a12696,a12698,a12700,a12702,a12704,a12706,a12708,a12710,a12712,a12714,a12716,a12718,a12720,
a12722,a12724,a12726,a12728,a12730,a12732,a12734,a12736,a12738,a12740,a12742,a12744,a12746,a12748,a12750,
a12752,a12754,a12756,a12758,a12760,a12762,a12764,a12766,a12768,a12770,a12772,a12774,a12776,a12778,a12780,
a12782,a12784,a12786,a12788,a12790,a12792,a12794,a12796,a12798,a12800,a12802,a12804,a12806,a12808,a12810,
a12812,a12814,a12816,a12818,a12820,a12822,a12824,a12826,a12828,a12830,a12832,a12834,a12836,a12838,a12840,
a12842,a12844,a12846,a12848,a12850,a12852,a12854,a12856,a12858,a12860,a12862,a12864,a12866,a12868,a12870,
a12872,a12874,a12876,a12878,a12880,a12882,a12884,a12886,a12888,a12890,a12892,a12894,a12896,a12898,a12900,
a12902,a12904,a12906,a12908,a12910,a12912,a12914,a12916,a12918,a12920,a12922,a12924,a12926,a12928,a12930,
a12932,a12934,a12936,a12938,a12940,a12942,a12944,a12946,a12948,a12950,a12952,a12954,a12956,a12958,a12960,
a12962,a12964,a12966,a12968,a12970,a12972,a12974,a12976,a12978,a12980,a12982,a12984,a12986,a12988,a12990,
a12992,a12994,a12996,a12998,a13000,a13002,a13004,a13006,a13008,a13010,a13012,a13014,a13016,a13018,a13020,
a13022,a13024,a13026,a13028,a13030,a13032,a13034,a13036,a13038,a13040,a13042,a13044,a13046,a13048,a13050,
a13052,a13054,a13056,a13058,a13060,a13062,a13064,a13066,a13068,a13070,a13072,a13074,a13076,a13078,a13080,
a13082,a13084,a13086,a13088,a13090,a13092,a13094,a13096,a13098,a13100,a13102,a13104,a13106,a13108,a13110,
a13112,a13114,a13116,a13118,a13120,a13122,a13124,a13126,a13128,a13130,a13132,a13134,a13136,a13138,a13140,
a13142,a13144,a13146,a13148,a13150,a13152,a13154,a13156,a13158,a13160,a13162,a13164,a13166,a13168,a13170,
a13172,a13174,a13176,a13178,a13180,a13182,a13184,a13186,a13188,a13190,a13192,a13194,a13196,a13198,a13200,
a13202,a13204,a13206,a13208,a13210,a13212,a13214,a13216,a13218,a13220,a13222,a13224,a13226,a13228,a13230,
a13232,a13234,a13236,a13238,a13240,a13242,a13244,a13246,a13248,a13250,a13252,a13254,a13256,a13258,a13260,
a13262,a13264,a13266,a13268,a13270,a13272,a13274,a13276,a13278,a13280,a13282,a13284,a13286,a13288,a13290,
a13292,a13294,a13296,a13298,a13300,a13302,a13304,a13306,a13308,a13310,a13312,a13314,a13316,a13318,a13320,
a13322,a13324,a13326,a13328,a13330,a13332,a13334,a13336,a13338,a13340,a13342,a13344,a13346,a13348,a13350,
a13352,a13354,a13356,a13358,a13360,a13362,a13364,a13366,a13368,a13370,a13372,a13374,a13376,a13378,a13380,
a13382,a13384,a13386,a13388,a13390,a13392,a13394,a13396,a13398,a13400,a13402,a13404,a13406,a13408,a13410,
a13412,a13414,a13416,a13418,a13420,a13422,a13424,a13426,a13428,a13430,a13432,a13434,a13436,a13438,a13440,
a13442,a13444,a13446,a13448,a13450,a13452,a13454,a13456,a13458,a13460,a13462,a13464,a13466,a13468,a13470,
a13472,a13474,a13476,a13478,a13480,a13482,a13484,a13486,a13488,a13490,a13492,a13494,a13496,a13498,a13500,
a13502,a13504,a13506,a13508,a13510,a13512,a13514,a13516,a13518,a13520,a13522,a13524,a13526,a13528,a13530,
a13532,a13534,a13536,a13538,a13540,a13542,a13544,a13546,a13548,a13550,a13552,a13554,a13556,a13558,a13560,
a13562,a13564,a13566,a13568,a13570,a13572,a13574,a13576,a13578,a13580,a13582,a13584,a13586,a13588,a13590,
a13592,a13594,a13596,a13598,a13600,a13602,a13604,a13606,a13608,a13610,a13612,a13614,a13616,a13618,a13620,
a13622,a13624,a13626,a13628,a13630,a13632,a13634,a13636,a13638,a13640,a13642,a13644,a13646,a13648,a13650,
a13652,a13654,a13656,a13658,a13660,a13662,a13664,a13666,a13668,a13670,a13672,a13674,a13676,a13678,a13680,
a13682,a13684,a13686,a13688,a13690,a13692,a13694,a13696,a13698,a13700,a13702,a13704,a13706,a13708,a13710,
a13712,a13714,a13716,a13718,a13720,a13722,a13724,a13726,a13728,a13730,a13732,a13734,a13736,a13738,a13740,
a13742,a13744,a13746,a13748,a13750,a13752,a13754,a13756,a13758,a13760,a13762,a13764,a13766,a13768,a13770,
a13772,a13774,a13776,a13778,a13780,a13782,a13784,a13786,a13788,a13790,a13792,a13794,a13796,a13798,a13800,
a13802,a13804,a13806,a13808,a13810,a13812,a13814,a13816,a13818,a13820,a13822,a13824,a13826,a13828,a13830,
a13832,a13834,a13836,a13838,a13840,a13842,a13844,a13846,a13848,a13850,a13852,a13854,a13856,a13858,a13860,
a13862,a13864,a13866,a13868,a13870,a13872,a13874,a13876,a13878,a13880,a13882,a13884,a13886,a13888,a13890,
a13892,a13894,a13896,a13898,a13900,a13902,a13904,a13906,a13908,a13910,a13912,a13914,a13916,a13918,a13920,
a13922,a13924,a13926,a13928,a13930,a13932,a13934,a13936,a13938,a13940,a13942,a13944,a13946,a13948,a13950,
a13952,a13954,a13956,a13958,a13960,a13962,a13964,a13966,a13968,a13970,a13972,a13974,a13976,a13978,a13980,
a13982,a13984,a13986,a13988,a13990,a13992,a13994,a13996,a13998,a14000,a14002,a14004,a14006,a14008,a14010,
a14012,a14014,a14016,a14018,a14020,a14022,a14024,a14026,a14028,a14030,a14032,a14034,a14036,a14038,a14040,
a14042,a14044,a14046,a14048,a14050,a14052,a14054,a14056,a14058,a14060,a14062,a14064,a14066,a14068,a14070,
a14072,a14074,a14076,a14078,a14080,a14082,a14084,a14086,a14088,a14090,a14092,a14094,a14096,a14098,a14100,
a14102,a14104,a14106,a14108,a14110,a14112,a14114,a14116,a14118,a14120,a14122,a14124,a14126,a14128,a14130,
a14132,a14134,a14136,a14138,a14140,a14142,a14144,a14146,a14148,a14150,a14152,a14154,a14156,a14158,a14160,
a14162,a14164,a14166,a14168,a14170,a14172,a14174,a14176,a14178,a14180,a14182,a14184,a14186,a14188,a14190,
a14192,a14194,a14196,a14198,a14200,a14202,a14204,a14206,a14208,a14210,a14212,a14214,a14216,a14218,a14220,
a14222,a14224,a14226,a14228,a14230,a14232,a14234,a14236,a14238,a14240,a14242,a14244,a14246,a14248,a14250,
a14252,a14254,a14256,a14258,a14260,a14262,a14264,a14266,a14268,a14270,a14272,a14274,a14276,a14278,a14280,
a14282,a14284,a14286,a14288,a14290,a14292,a14294,a14296,a14298,a14300,a14302,a14304,a14306,a14308,a14310,
a14312,a14314,a14316,a14318,a14320,a14322,a14324,a14326,a14328,a14330,a14332,a14334,a14336,a14338,a14340,
a14342,a14344,a14346,a14348,a14350,a14352,a14354,a14356,a14358,a14360,a14362,a14364,a14366,a14368,a14370,
a14372,a14374,a14376,a14378,a14380,a14382,a14384,a14386,a14388,a14390,a14392,a14394,a14396,a14398,a14400,
a14402,a14404,a14406,a14408,a14410,a14412,a14414,a14416,a14418,a14420,a14422,a14424,a14426,a14428,a14430,
a14432,a14434,a14436,a14438,a14440,a14442,a14444,a14446,a14448,a14450,a14452,a14454,a14456,a14458,a14460,
a14462,a14464,a14466,a14468,a14470,a14472,a14474,a14476,a14478,a14480,a14482,a14484,a14486,a14488,a14490,
a14492,a14494,a14496,a14498,a14500,a14502,a14504,a14506,a14508,a14510,a14512,a14514,a14516,a14518,a14520,
a14522,a14524,a14526,a14528,a14530,a14532,a14534,a14536,a14538,a14540,a14542,a14544,a14546,a14548,a14550,
a14552,a14554,a14556,a14558,a14560,a14562,a14564,a14566,a14568,a14570,a14572,a14574,a14576,a14578,a14580,
a14582,a14584,a14586,a14588,a14590,a14592,a14594,a14596,a14598,a14600,a14602,a14604,a14606,a14608,a14610,
a14612,a14614,a14616,a14618,a14620,a14622,a14624,a14626,a14628,a14630,a14632,a14634,a14636,a14638,a14640,
a14642,a14644,a14646,a14648,a14650,a14652,a14654,a14656,a14658,a14660,a14662,a14664,a14666,a14668,a14670,
a14672,a14674,a14676,a14678,a14680,a14682,a14684,a14686,a14688,a14690,a14692,a14694,a14696,a14698,a14700,
a14702,a14704,a14706,a14708,a14710,a14712,a14714,a14716,a14718,a14720,a14722,a14724,a14726,a14728,a14730,
a14732,a14734,a14736,a14738,a14740,a14742,a14744,a14746,a14748,a14750,a14752,a14754,a14756,a14758,a14760,
a14762,a14764,a14766,a14768,a14770,a14772,a14774,a14776,a14778,a14780,a14782,a14784,a14786,a14788,a14790,
a14792,a14794,a14796,a14798,a14800,a14802,a14804,a14806,a14808,a14810,a14812,a14814,a14816,a14818,a14820,
a14822,a14824,a14826,a14828,a14830,a14832,a14834,a14836,a14838,a14840,a14842,a14844,a14846,a14848,a14850,
a14852,a14854,a14856,a14858,a14860,a14862,a14864,a14866,a14868,a14870,a14872,a14874,a14876,a14878,a14880,
a14882,a14884,a14886,a14888,a14890,a14892,a14894,a14896,a14898,a14900,a14902,a14904,a14906,a14908,a14910,
a14912,a14914,a14916,a14918,a14920,a14922,a14924,a14926,a14928,a14930,a14932,a14934,a14936,a14938,a14940,
a14942,a14944,a14946,a14948,a14950,a14952,a14954,a14956,a14958,a14960,a14962,a14964,a14966,a14968,a14970,
a14972,a14974,a14976,a14978,a14980,a14982,a14984,a14986,a14988,a14990,a14992,a14994,a14996,a14998,a15000,
a15002,a15004,a15006,a15008,a15010,a15012,a15014,a15016,a15018,a15020,a15022,a15024,a15026,a15028,a15030,
a15032,a15034,a15036,a15038,a15040,a15042,a15044,a15046,a15048,a15050,a15052,a15054,a15056,a15058,a15060,
a15062,a15064,a15066,a15068,a15070,a15072,a15074,a15076,a15078,a15080,a15082,a15084,a15086,a15088,a15090,
a15092,a15094,a15096,a15098,a15100,a15102,a15104,a15106,a15108,a15110,a15112,a15114,a15116,a15118,a15120,
a15122,a15124,a15126,a15128,a15130,a15132,a15134,a15136,a15138,a15140,a15142,a15144,a15146,a15148,a15150,
a15152,a15154,a15156,a15158,a15160,a15162,a15164,a15166,a15168,a15170,a15172,a15174,a15176,a15178,a15180,
a15182,a15184,a15186,a15188,a15190,a15192,a15194,a15196,a15198,a15200,a15202,a15204,a15206,a15208,a15210,
a15212,a15214,a15216,a15218,a15220,a15222,a15224,a15226,a15228,a15230,a15232,a15234,a15236,a15238,a15240,
a15242,a15244,a15246,a15248,a15250,a15252,a15254,a15256,a15258,a15260,a15262,a15264,a15266,a15268,a15270,
a15272,a15274,a15276,a15278,a15280,a15282,a15284,a15286,a15288,a15290,a15292,a15294,a15296,a15298,a15300,
a15302,a15304,a15306,a15308,a15310,a15312,a15314,a15316,a15318,a15320,a15322,a15324,a15326,a15328,a15330,
a15332,a15334,a15336,a15338,a15340,a15342,a15344,a15346,a15348,a15350,a15352,a15354,a15356,a15358,a15360,
a15362,a15364,a15366,a15368,a15370,a15372,a15374,a15376,a15378,a15380,a15382,a15384,a15386,a15388,a15390,
a15392,a15394,a15396,a15398,a15400,a15402,a15404,a15406,a15408,a15410,a15412,a15414,a15416,a15418,a15420,
a15422,a15424,a15426,a15428,a15430,a15432,a15434,a15436,a15438,a15440,a15442,a15444,a15446,a15448,a15450,
a15452,a15454,a15456,a15458,a15460,a15462,a15464,a15466,a15468,a15470,a15472,a15474,a15476,a15478,a15480,
a15482,a15484,a15486,a15488,a15490,a15492,a15494,a15496,a15498,a15500,a15502,a15504,a15506,a15508,a15510,
a15512,a15514,a15516,a15518,a15520,a15522,a15524,a15526,a15528,a15530,a15532,a15534,a15536,a15538,a15540,
a15542,a15544,a15546,a15548,a15550,a15552,a15554,a15556,a15558,a15560,a15562,a15564,a15566,a15568,a15570,
a15572,a15574,a15576,a15578,a15580,a15582,a15584,a15586,a15588,a15590,a15592,a15594,a15596,a15598,a15600,
a15602,a15604,a15606,a15608,a15610,a15612,a15614,a15616,a15618,a15620,a15622,a15624,a15626,a15628,a15630,
a15632,a15634,a15636,a15638,a15640,a15642,a15644,a15646,a15648,a15650,a15652,a15654,a15656,a15658,a15660,
a15662,a15664,a15666,a15668,a15670,a15672,a15674,a15676,a15678,a15680,a15682,a15684,a15686,a15688,a15690,
a15692,a15694,a15696,a15698,a15700,a15702,a15704,a15706,a15708,a15710,a15712,a15714,a15716,a15718,a15720,
a15722,a15724,a15726,a15728,a15730,a15732,a15734,a15736,a15738,a15740,a15742,a15744,a15746,a15748,a15750,
a15752,a15754,a15756,a15758,a15760,a15762,a15764,a15766,a15768,a15770,a15772,a15774,a15776,a15778,a15780,
a15782,a15784,a15786,a15788,a15790,a15792,a15794,a15796,a15798,a15800,a15802,a15804,a15806,a15808,a15810,
a15812,a15814,a15816,a15818,a15820,a15822,a15824,a15826,a15828,a15830,a15832,a15834,a15836,a15838,a15840,
a15842,a15844,a15846,a15848,a15850,a15852,a15854,a15856,a15858,a15860,a15862,a15864,a15866,a15868,a15870,
a15872,a15874,a15876,a15878,a15880,a15882,a15884,a15886,a15888,a15890,a15892,a15894,a15896,a15898,a15900,
a15902,a15904,a15906,a15908,a15910,a15912,a15914,a15916,a15918,a15920,a15922,a15924,a15926,a15928,a15930,
a15932,a15934,a15936,a15938,a15940,a15942,a15944,a15946,a15948,a15950,a15952,a15954,a15956,a15958,a15960,
a15962,a15964,a15966,a15968,a15970,a15972,a15974,a15976,a15978,a15980,a15982,a15984,a15986,a15988,a15990,
a15992,a15994,a15996,a15998,a16000,a16002,a16004,a16006,a16008,a16010,a16012,a16014,a16016,a16018,a16020,
a16022,a16024,a16026,a16028,a16030,a16032,a16034,a16036,a16038,a16040,a16042,a16044,a16046,a16048,a16050,
a16052,a16054,a16056,a16058,a16060,a16062,a16064,a16066,a16068,a16070,a16072,a16074,a16076,a16078,a16080,
a16082,a16084,a16086,a16088,a16090,a16092,a16094,a16096,a16098,a16100,a16102,a16104,a16106,a16108,a16110,
a16112,a16114,a16116,a16118,a16120,a16122,a16124,a16126,a16128,a16130,a16132,a16134,a16136,a16138,a16140,
a16142,a16144,a16146,a16148,a16150,a16152,a16154,a16156,a16158,a16160,a16162,a16164,a16166,a16168,a16170,
a16172,a16174,a16176,a16178,a16180,a16182,a16184,a16186,a16188,a16190,a16192,a16194,a16196,a16198,a16200,
a16202,a16204,a16206,a16208,a16210,a16212,a16214,a16216,a16218,a16220,a16222,a16224,a16226,a16228,a16230,
a16232,a16234,a16236,a16238,a16240,a16242,a16244,a16246,a16248,a16250,a16252,a16254,a16256,a16258,a16260,
a16262,a16264,a16266,a16268,a16270,a16272,a16274,a16276,a16278,a16280,a16282,a16284,a16286,a16288,a16290,
a16292,a16294,a16296,a16298,a16300,a16302,a16304,a16306,a16308,a16310,a16312,a16314,a16316,a16318,a16320,
a16322,a16324,a16326,a16328,a16330,a16332,a16334,a16336,a16338,a16340,a16342,a16344,a16346,a16348,a16350,
a16352,a16354,a16356,a16358,a16360,a16362,a16364,a16366,a16368,a16370,a16372,a16374,a16376,a16378,a16380,
a16382,a16384,a16386,a16388,a16390,a16392,a16394,a16396,a16398,a16400,a16402,a16404,a16406,a16408,a16410,
a16412,a16414,a16416,a16418,a16420,a16422,a16424,a16426,a16428,a16430,a16432,a16434,a16436,a16438,a16440,
a16442,a16444,a16446,a16448,a16450,a16452,a16454,a16456,a16458,a16460,a16462,a16464,a16466,a16468,a16470,
a16472,a16474,a16476,a16478,a16480,a16482,a16484,a16486,a16488,a16490,a16492,a16494,a16496,a16498,a16500,
a16502,a16504,a16506,a16508,a16510,a16512,a16514,a16516,a16518,a16520,a16522,a16524,a16526,a16528,a16530,
a16532,a16534,a16536,a16538,a16540,a16542,a16544,a16546,a16548,a16550,a16552,a16554,a16556,a16558,a16560,
a16562,a16564,a16566,a16568,a16570,a16572,a16574,a16576,a16578,a16580,a16582,a16584,a16586,a16588,a16590,
a16592,a16594,a16596,a16598,a16600,a16602,a16604,a16606,a16608,a16610,a16612,a16614,a16616,a16618,a16620,
a16622,a16624,a16626,a16628,a16630,a16632,a16634,a16636,a16638,a16640,a16642,a16644,a16646,a16648,a16650,
a16652,a16654,a16656,a16658,a16660,a16662,a16664,a16666,a16668,a16670,a16672,a16674,a16676,a16678,a16680,
a16682,a16684,a16686,a16688,a16690,a16692,a16694,a16696,a16698,a16700,a16702,a16704,a16706,a16708,a16710,
a16712,a16714,a16716,a16718,a16720,a16722,a16724,a16726,a16728,a16730,a16732,a16734,a16736,a16738,a16740,
a16742,a16744,a16746,a16748,a16750,a16752,a16754,a16756,a16758,a16760,a16762,a16764,a16766,a16768,a16770,
a16772,a16774,a16776,a16778,a16780,a16782,a16784,a16786,a16788,a16790,a16792,a16794,a16796,a16798,a16800,
a16802,a16804,a16806,a16808,a16810,a16812,a16814,a16816,a16818,a16820,a16822,a16824,a16826,a16828,a16830,
a16832,a16834,a16836,a16838,a16840,a16842,a16844,a16846,a16848,a16850,a16852,a16854,a16856,a16858,a16860,
a16862,a16864,a16866,a16868,a16870,a16872,a16874,a16876,a16878,a16880,a16882,a16884,a16886,a16888,a16890,
a16892,a16894,a16896,a16898,a16900,a16902,a16904,a16906,a16908,a16910,a16912,a16914,a16916,a16918,a16920,
a16922,a16924,a16926,a16928,a16930,a16932,a16934,a16936,a16938,a16940,a16942,a16944,a16946,a16948,a16950,
a16952,a16954,a16956,a16958,a16960,a16962,a16964,a16966,a16968,a16970,a16972,a16974,a16976,a16978,a16980,
a16982,a16984,a16986,a16988,a16990,a16992,a16994,a16996,a16998,a17000,a17002,a17004,a17006,a17008,a17010,
a17012,a17014,a17016,a17018,a17020,a17022,a17024,a17026,a17028,a17030,a17032,a17034,a17036,a17038,a17040,
a17042,a17044,a17046,a17048,a17050,a17052,a17054,a17056,a17058,a17060,a17062,a17064,a17066,a17068,a17070,
a17072,a17074,a17076,a17078,a17080,a17082,a17084,a17086,a17088,a17090,a17092,a17094,a17096,a17098,a17100,
a17102,a17104,a17106,a17108,a17110,a17112,a17114,a17116,a17118,a17120,a17122,a17124,a17126,a17128,a17130,
a17132,a17134,a17136,a17138,a17140,a17142,a17144,a17146,a17148,a17150,a17152,a17154,a17156,a17158,a17160,
a17162,a17164,a17166,a17168,a17170,a17172,a17174,a17176,a17178,a17180,a17182,a17184,a17186,a17188,a17190,
a17192,a17194,a17196,a17198,a17200,a17202,a17204,a17206,a17208,a17210,a17212,a17214,a17216,a17218,a17220,
a17222,a17224,a17226,a17228,a17230,a17232,a17234,a17236,a17238,a17240,a17242,a17244,a17246,a17248,a17250,
a17252,a17254,a17256,a17258,a17260,a17262,a17264,a17266,a17268,a17270,a17272,a17274,a17276,a17278,a17280,
a17282,a17284,a17286,a17288,a17290,a17292,a17294,a17296,a17298,a17300,a17302,a17304,a17306,a17308,a17310,
a17312,a17314,a17316,a17318,a17320,a17322,a17324,a17326,a17328,a17330,a17332,a17334,a17336,a17338,a17340,
a17342,a17344,a17346,a17348,a17350,a17352,a17354,a17356,a17358,a17360,a17362,a17364,a17366,a17368,a17370,
a17372,a17374,a17376,a17378,a17380,a17382,a17384,a17386,a17388,a17390,a17392,a17394,a17396,a17398,a17400,
a17402,a17404,a17406,a17408,a17410,a17412,a17414,a17416,a17418,a17420,a17422,a17424,a17426,a17428,a17430,
a17432,a17434,a17436,a17438,a17440,a17442,a17444,a17446,a17448,a17450,a17452,a17454,a17456,a17458,a17460,
a17462,a17464,a17466,a17468,a17470,a17472,a17474,a17476,a17478,a17480,a17482,a17484,a17486,a17488,a17490,
a17492,a17494,a17496,a17498,a17500,a17502,a17504,a17506,a17508,a17510,a17512,a17514,a17516,a17518,a17520,
a17522,a17524,a17526,a17528,a17530,a17532,a17534,a17536,a17538,a17540,a17542,a17544,a17546,a17548,a17550,
a17552,a17554,a17556,a17558,a17560,a17562,a17564,a17566,a17568,a17570,a17572,a17574,a17576,a17578,a17580,
a17582,a17584,a17586,a17588,a17590,a17592,a17594,a17596,a17598,a17600,a17602,a17604,a17606,a17608,a17610,
a17612,a17614,a17616,a17618,a17620,a17622,a17624,a17626,a17628,a17630,a17632,a17634,a17636,a17638,a17640,
a17642,a17644,a17646,a17648,a17650,a17652,a17654,a17656,a17658,a17660,a17662,a17664,a17666,a17668,a17670,
a17672,a17674,a17676,a17678,a17680,a17682,a17684,a17686,a17688,a17690,a17692,a17694,a17696,a17698,a17700,
a17702,a17704,a17706,a17708,a17710,a17712,a17714,a17716,a17718,a17720,a17722,a17724,a17726,a17728,a17730,
a17732,a17734,a17736,a17738,a17740,a17742,a17744,a17746,a17748,a17750,a17752,a17754,a17756,a17758,a17760,
a17762,a17764,a17766,a17768,a17770,a17772,a17774,a17776,a17778,a17780,a17782,a17784,a17786,a17788,a17790,
a17792,a17794,a17796,a17798,a17800,a17802,a17804,a17806,a17808,a17810,a17812,a17814,a17816,a17818,a17820,
a17822,a17824,a17826,a17828,a17830,a17832,a17834,a17836,a17838,a17840,a17842,a17844,a17846,a17848,a17850,
a17852,a17854,a17856,a17858,a17860,a17862,a17864,a17866,a17868,a17870,a17872,a17874,a17876,a17878,a17880,
a17882,a17884,a17886,a17888,a17890,a17892,a17894,a17896,a17898,a17900,a17902,a17904,a17906,a17908,a17910,
a17912,a17914,a17916,a17918,a17920,a17922,a17924,a17926,a17928,a17930,a17932,a17934,a17936,a17938,a17940,
a17942,a17944,a17946,a17948,a17950,a17952,a17954,a17956,a17958,a17960,a17962,a17964,a17966,a17968,a17970,
a17972,a17974,a17976,a17978,a17980,a17982,a17984,a17986,a17988,a17990,a17992,a17994,a17996,a17998,a18000,
a18002,a18004,a18006,a18008,a18010,a18012,a18014,a18016,a18018,a18020,a18022,a18024,a18026,a18028,a18030,
a18032,a18034,a18036,a18038,a18040,a18042,a18044,a18046,a18048,a18050,a18052,a18054,a18056,a18058,a18060,
a18062,a18064,a18066,a18068,a18070,a18072,a18074,a18076,a18078,a18080,a18082,a18084,a18086,a18088,a18090,
a18092,a18094,a18096,a18098,a18100,a18102,a18104,a18106,a18108,a18110,a18112,a18114,a18116,a18118,a18120,
a18122,a18124,a18126,a18128,a18130,a18132,a18134,a18136,a18138,a18140,a18142,a18144,a18146,a18148,a18150,
a18152,a18154,a18156,a18158,a18160,a18162,a18164,a18166,a18168,a18170,a18172,a18174,a18176,a18178,a18180,
a18182,a18184,a18186,a18188,a18190,a18192,a18194,a18196,a18198,a18200,a18202,a18204,a18206,a18208,a18210,
a18212,a18214,a18216,a18218,a18220,a18222,a18224,a18226,a18228,a18230,a18232,a18234,a18236,a18238,a18240,
a18242,a18244,a18246,a18248,a18250,a18252,a18254,a18256,a18258,a18260,a18262,a18264,a18266,a18268,a18270,
a18272,a18274,a18276,a18278,a18280,a18282,a18284,a18286,a18288,a18290,a18292,a18294,a18296,a18298,a18300,
a18302,a18304,a18306,a18308,a18310,a18312,a18314,a18316,a18318,a18320,a18322,a18324,a18326,a18328,a18330,
a18332,a18334,a18336,a18338,a18340,a18342,a18344,a18346,a18348,a18350,a18352,a18354,a18356,a18358,a18360,
a18362,a18364,a18366,a18368,a18370,a18372,a18374,a18376,a18378,a18380,a18382,a18384,a18386,a18388,a18390,
a18392,a18394,a18396,a18398,a18400,a18402,a18404,a18406,a18408,a18410,a18412,a18414,a18416,a18418,a18420,
a18422,a18424,a18426,a18428,a18430,a18432,a18434,a18436,a18438,a18440,a18442,a18444,a18446,a18448,a18450,
a18452,a18454,a18456,a18458,a18460,a18462,a18464,a18466,a18468,a18470,a18472,a18474,a18476,a18478,a18480,
a18482,a18484,a18486,a18488,a18490,a18492,a18494,a18496,a18498,a18500,a18502,a18504,a18506,a18508,a18510,
a18512,a18514,a18516,a18518,a18520,a18522,a18524,a18526,a18528,a18530,a18532,a18534,a18536,a18538,a18540,
a18542,a18544,a18546,a18548,a18550,a18552,a18554,a18556,a18558,a18560,a18562,a18564,a18566,a18568,a18570,
a18572,a18574,a18576,a18578,a18580,a18582,a18584,a18586,a18588,a18590,a18592,a18594,a18596,a18598,a18600,
a18602,a18604,a18606,a18608,a18610,a18612,a18614,a18616,a18618,a18620,a18622,a18624,a18626,a18628,a18630,
a18632,a18634,a18636,a18638,a18640,a18642,a18644,a18646,a18648,a18650,a18652,a18654,a18656,a18658,a18660,
a18662,a18664,a18666,a18668,a18670,a18672,a18674,a18676,a18678,a18680,a18682,a18684,a18686,a18688,a18690,
a18692,a18694,a18696,a18698,a18700,a18702,a18704,a18706,a18708,a18710,a18712,a18714,a18716,a18718,a18720,
a18722,a18724,a18726,a18728,a18730,a18732,a18734,a18736,a18738,a18740,a18742,a18744,a18746,a18748,a18750,
a18752,a18754,a18756,a18758,a18760,a18762,a18764,a18766,a18768,a18770,a18772,a18774,a18776,a18778,a18780,
a18782,a18784,a18786,a18788,a18790,a18792,a18794,a18796,a18798,a18800,a18802,a18804,a18806,a18808,a18810,
a18812,a18814,a18816,a18818,a18820,a18822,a18824,a18826,a18828,a18830,a18832,a18834,a18836,a18838,a18840,
a18842,a18844,a18846,a18848,a18850,a18852,a18854,a18856,a18858,a18860,a18862,a18864,a18866,a18868,a18870,
a18872,a18874,a18876,a18878,a18880,a18882,a18884,a18886,a18888,a18890,a18892,a18894,a18896,a18898,a18900,
a18902,a18904,a18906,a18908,a18910,a18912,a18914,a18916,a18918,a18920,a18922,a18924,a18926,a18928,a18930,
a18932,a18934,a18936,a18938,a18940,a18942,a18944,a18946,a18948,a18950,a18952,a18954,a18956,a18958,a18960,
a18962,a18964,a18966,a18968,a18970,a18972,a18974,a18976,a18978,a18980,a18982,a18984,a18986,a18988,a18990,
a18992,a18994,a18996,a18998,a19000,a19002,a19004,a19006,a19008,a19010,a19012,a19014,a19016,a19018,a19020,
a19022,a19024,a19026,a19028,a19030,a19032,a19034,a19036,a19038,a19040,a19042,a19044,a19046,a19048,a19050,
a19052,a19054,a19056,a19058,a19060,a19062,a19064,a19066,a19068,a19070,a19072,a19074,a19076,a19078,a19080,
a19082,a19084,a19086,a19088,a19090,a19092,a19094,a19096,a19098,a19100,a19102,a19104,a19106,a19108,a19110,
a19112,a19114,a19116,a19118,a19120,a19122,a19124,a19126,a19128,a19130,a19132,a19134,a19136,a19138,a19140,
a19142,a19144,a19146,a19148,a19150,a19152,a19154,a19156,a19158,a19160,a19162,a19164,a19166,a19168,a19170,
a19172,a19174,a19176,a19178,a19180,a19182,a19184,a19186,a19188,a19190,a19192,a19194,a19196,a19198,a19200,
a19202,a19204,a19206,a19208,a19210,a19212,a19214,a19216,a19218,a19220,a19222,a19224,a19226,a19228,a19230,
a19232,a19234,a19236,a19238,a19240,a19242,a19244,a19246,a19248,a19250,a19252,a19254,a19256,a19258,a19260,
a19262,a19264,a19266,a19268,a19270,a19272,a19274,a19276,a19278,a19280,a19282,a19284,a19286,a19288,a19290,
a19292,a19294,a19296,a19298,a19300,a19302,a19304,a19306,a19308,a19310,a19312,a19314,a19316,a19318,a19320,
a19322,a19324,a19326,a19328,a19330,a19332,a19334,a19336,a19338,a19340,a19342,a19344,a19346,a19348,a19350,
a19352,a19354,a19356,a19358,a19360,a19362,a19364,a19366,a19368,a19370,a19372,a19374,a19376,a19378,a19380,
a19382,a19384,a19386,a19388,a19390,a19392,a19394,a19396,a19398,a19400,a19402,a19404,a19406,a19408,a19410,
a19412,a19414,a19416,a19418,a19420,a19422,a19424,a19426,a19428,a19430,a19432,a19434,a19436,a19438,a19440,
a19442,a19444,a19446,a19448,a19450,a19452,a19454,a19456,a19458,a19460,a19462,a19464,a19466,a19468,a19470,
a19474,a19476,a19478,a19480,a19482,a19484,a19486,a19488,a19490,a19492,a19494,a19496,a19498,a19500,a19502,
a19504,a19506,a19508,a19510,a19512,a19514,a19516,a19518,a19520,a19522,a19524,a19526,a19528,a19530,a19532,
a19534,a19536,a19538,a19540,a19542,a19544,a19546,a19548,a19550,a19552,a19554,a19556,a19558,a19560,a19562,
a19564,a19566,a19568,a19570,a19572,a19574,a19576,a19578,a19580,a19582,a19584,a19586,a19588,a19590,a19592,
a19594,a19596,a19598,a19600,a19602,a19604,a19606,a19608,a19610,a19612,a19614,a19616,a19618,a19620,a19622,
a19624,a19626,a19628,a19630,a19632,a19634,a19636,a19638,a19640,a19642,a19644,a19646,a19648,a19650,a19652,
a19654,a19656,a19658,a19660,a19662,a19664,a19666,a19668,a19670,a19672,a19674,a19676,a19678,a19680,a19682,
a19684,a19686,a19688,a19690,a19692,a19694,a19696,a19698,a19700,a19702,a19704,a19706,a19708,a19710,a19712,
a19714,a19716,a19718,a19720,a19722,a19724,a19726,a19728,a19730,a19732,a19734,a19736,a19738,a19740,a19742,
a19744,a19746,a19748,a19750,a19752,a19754,a19756,a19758,a19760,a19762,a19764,a19766,a19768,a19770,a19772,
a19774,a19776,a19778,a19780,a19782,a19784,a19786,a19788,a19790,a19792,a19794,a19796,a19798,a19800,a19802,
a19804,a19806,a19808,a19810,a19812,a19814,a19816,a19818,a19820,a19822,a19824,a19826,a19828,a19830,a19832,
a19834,a19836,a19838,a19840,a19842,a19844,a19846,a19848,a19850,a19852,a19854,a19856,a19858,a19860,a19862,
a19864,a19866,a19868,a19870,a19872,a19874,a19876,a19878,a19880,a19882,a19884,a19886,a19888,a19890,a19892,
a19894,a19896,a19898,a19900,a19902,a19904,a19906,a19908,a19910,a19912,a19914,a19916,a19918,a19920,a19922,
a19924,a19926,a19928,a19930,a19932,a19934,a19936,a19938,a19940,a19942,a19944,a19946,a19948,a19950,a19952,
a19954,a19956,a19958,a19960,a19962,a19964,a19966,a19968,a19970,a19972,a19974,a19976,a19978,a19980,a19982,
a19984,a19986,a19988,a19990,a19992,a19994,a19996,a19998,a20000,a20002,a20004,a20006,a20008,a20010,a20012,
a20014,a20016,a20018,a20020,a20022,a20024,a20026,a20028,a20030,a20032,a20034,a20036,a20038,a20040,a20042,
a20044,a20046,a20048,a20050,a20052,a20054,a20056,a20058,a20060,a20062,a20064,a20066,a20068,a20070,a20072,
a20074,a20076,a20078,a20080,a20082,a20084,a20086,a20088,a20090,a20092,a20094,a20096,a20098,a20100,a20102,
a20104,a20106,a20108,a20110,a20112,a20114,a20116,a20118,a20120,a20122,a20124,a20126,a20128,a20130,a20132,
a20134,a20136,a20138,a20140,a20142,a20144,a20146,a20148,a20150,a20152,a20154,a20156,a20158,a20160,a20162,
a20164,a20166,a20168,a20170,a20172,a20174,a20176,a20178,a20180,a20182,a20184,a20186,a20188,a20190,a20192,
a20194,a20196,a20198,a20200,a20202,a20204,a20206,a20208,a20210,a20212,a20214,a20216,a20218,a20220,a20222,
a20224,a20226,a20228,a20230,a20232,a20234,a20236,a20238,a20240,a20242,a20244,a20246,a20248,a20250,a20252,
a20254,a20256,a20258,a20260,a20262,a20264,a20266,a20268,a20270,a20272,a20274,a20276,a20278,a20280,a20282,
a20284,a20286,a20288,a20290,a20292,a20294,a20296,a20298,a20300,a20302,a20304,a20306,a20308,a20310,a20312,
a20314,a20316,a20318,a20320,a20322,a20324,a20326,a20328,a20330,a20332,a20334,a20336,a20338,a20340,a20342,
a20344,a20346,a20348,a20350,a20352,a20354,a20356,p0,p1,p2,p3,p4;

reg l164,l166,l168,l170,l172,l174,l176,l178,l180,l182,l184,l186,l188,l190,l192,
l194,l196,l198,l200,l202,l204,l206,l208,l210,l212,l214,l216,l218,l220,l222,
l224,l226,l228,l230,l232,l234,l236,l238,l240,l242,l244,l246,l248,l250,l252,
l254,l256,l258,l260,l262,l264,l266,l268,l270,l272,l274,l276,l278,l280,l282,
l284,l286,l288,l290,l292,l294,l296,l298,l300,l302,l304,l306,l308,l310,l312,
l314,l316,l318,l320,l322,l324,l326,l328,l330,l332,l334,l336,l338,l340;

initial
begin
   l164 = 0;
   l166 = 0;
   l168 = 0;
   l170 = 0;
   l172 = 0;
   l174 = 1;
   l176 = 0;
   l178 = 1;
   l180 = 0;
   l182 = 0;
   l184 = 0;
   l186 = 0;
   l188 = 0;
   l190 = 0;
   l192 = 0;
   l194 = 0;
   l196 = 0;
   l198 = 0;
   l200 = 0;
   l202 = 0;
   l204 = 0;
   l206 = 0;
   l208 = 0;
   l210 = 0;
   l212 = 0;
   l214 = 0;
   l216 = 0;
   l218 = 0;
   l220 = 0;
   l222 = 0;
   l224 = 0;
   l226 = 0;
   l228 = 0;
   l230 = 0;
   l232 = 0;
   l234 = 0;
   l236 = 0;
   l238 = 0;
   l240 = 0;
   l242 = 0;
   l244 = 0;
   l246 = 0;
   l248 = 0;
   l250 = 0;
   l252 = 0;
   l254 = 0;
   l256 = 0;
   l258 = 0;
   l260 = 0;
   l262 = 0;
   l264 = 0;
   l266 = 0;
   l268 = 0;
   l270 = 0;
   l272 = 0;
   l274 = 0;
   l276 = 0;
   l278 = 0;
   l280 = 0;
   l282 = 0;
   l284 = 0;
   l286 = 0;
   l288 = 0;
   l290 = 0;
   l292 = 0;
   l294 = 0;
   l296 = 0;
   l298 = 0;
   l300 = 0;
   l302 = 0;
   l304 = 0;
   l306 = 0;
   l308 = 0;
   l310 = 0;
   l312 = 0;
   l314 = 0;
   l316 = 0;
   l318 = 0;
   l320 = 0;
   l322 = 2;
   l324 = 0;
   l326 = 0;
   l328 = 0;
   l330 = 0;
   l332 = 0;
   l334 = 0;
   l336 = 0;
   l338 = 0;
   l340 = 0;
end

always @(posedge i2)
   l164 <= i2;

always @(posedge i4)
   l166 <= i4;

always @(posedge i6)
   l168 <= i6;

always @(posedge i8)
   l170 <= i8;

always @(posedge i10)
   l172 <= i10;

always @(posedge na342)
   l174 <= na342;

always @(posedge a344)
   l176 <= a344;

always @(posedge na346)
   l178 <= na346;

always @(posedge a348)
   l180 <= a348;

always @(posedge a350)
   l182 <= a350;

always @(posedge i12)
   l184 <= i12;

always @(posedge i14)
   l186 <= i14;

always @(posedge i16)
   l188 <= i16;

always @(posedge i18)
   l190 <= i18;

always @(posedge i20)
   l192 <= i20;

always @(posedge i22)
   l194 <= i22;

always @(posedge i24)
   l196 <= i24;

always @(posedge i26)
   l198 <= i26;

always @(posedge i28)
   l200 <= i28;

always @(posedge i30)
   l202 <= i30;

always @(posedge i32)
   l204 <= i32;

always @(posedge i34)
   l206 <= i34;

always @(posedge i36)
   l208 <= i36;

always @(posedge i38)
   l210 <= i38;

always @(posedge i40)
   l212 <= i40;

always @(posedge i42)
   l214 <= i42;

always @(posedge i44)
   l216 <= i44;

always @(posedge i46)
   l218 <= i46;

always @(posedge i48)
   l220 <= i48;

always @(posedge i50)
   l222 <= i50;

always @(posedge i52)
   l224 <= i52;

always @(posedge i54)
   l226 <= i54;

always @(posedge i56)
   l228 <= i56;

always @(posedge i58)
   l230 <= i58;

always @(posedge i60)
   l232 <= i60;

always @(posedge i62)
   l234 <= i62;

always @(posedge i64)
   l236 <= i64;

always @(posedge i66)
   l238 <= i66;

always @(posedge i68)
   l240 <= i68;

always @(posedge i70)
   l242 <= i70;

always @(posedge i72)
   l244 <= i72;

always @(posedge i74)
   l246 <= i74;

always @(posedge i76)
   l248 <= i76;

always @(posedge i78)
   l250 <= i78;

always @(posedge i80)
   l252 <= i80;

always @(posedge i82)
   l254 <= i82;

always @(posedge i84)
   l256 <= i84;

always @(posedge i86)
   l258 <= i86;

always @(posedge i88)
   l260 <= i88;

always @(posedge i90)
   l262 <= i90;

always @(posedge i92)
   l264 <= i92;

always @(posedge i94)
   l266 <= i94;

always @(posedge i96)
   l268 <= i96;

always @(posedge i98)
   l270 <= i98;

always @(posedge i100)
   l272 <= i100;

always @(posedge i102)
   l274 <= i102;

always @(posedge i104)
   l276 <= i104;

always @(posedge i106)
   l278 <= i106;

always @(posedge i108)
   l280 <= i108;

always @(posedge i110)
   l282 <= i110;

always @(posedge i112)
   l284 <= i112;

always @(posedge i114)
   l286 <= i114;

always @(posedge i116)
   l288 <= i116;

always @(posedge i118)
   l290 <= i118;

always @(posedge i120)
   l292 <= i120;

always @(posedge i122)
   l294 <= i122;

always @(posedge i124)
   l296 <= i124;

always @(posedge i126)
   l298 <= i126;

always @(posedge i128)
   l300 <= i128;

always @(posedge i130)
   l302 <= i130;

always @(posedge i132)
   l304 <= i132;

always @(posedge i134)
   l306 <= i134;

always @(posedge i136)
   l308 <= i136;

always @(posedge i138)
   l310 <= i138;

always @(posedge i140)
   l312 <= i140;

always @(posedge i142)
   l314 <= i142;

always @(posedge i144)
   l316 <= i144;

always @(posedge i146)
   l318 <= i146;

always @(posedge i148)
   l320 <= i148;

always @(posedge z0)
   l322 <= z0;

always @(posedge i150)
   l324 <= i150;

always @(posedge i152)
   l326 <= i152;

always @(posedge i154)
   l328 <= i154;

always @(posedge i156)
   l330 <= i156;

always @(posedge i158)
   l332 <= i158;

always @(posedge i160)
   l334 <= i160;

always @(posedge i162)
   l336 <= i162;

always @(posedge a19472)
   l338 <= a19472;

always @(posedge c1)
   l340 <= c1;


assign na342 = ~a342;
assign a344 = l340 & l166;
assign na346 = ~a346;
assign a348 = l340 & l170;
assign a350 = l340 & l172;
assign z0 = l322;
assign a19472 = ~a19470 & ~a842;
assign c1 = 1;
assign a342 = l340 & ~l164;
assign a346 = l340 & ~l168;
assign a352 = i74 & ~i72;
assign a354 = a352 & ~i70;
assign a356 = ~i74 & ~i72;
assign a358 = a356 & i70;
assign a360 = ~a352 & ~i70;
assign a362 = ~a360 & ~a358;
assign a364 = a362 & ~a354;
assign a366 = ~a364 & ~i62;
assign a368 = a364 & i62;
assign a370 = ~a368 & ~a366;
assign a372 = i20 & i18;
assign a374 = a372 & ~i16;
assign a376 = a374 & ~i34;
assign a378 = ~a374 & i34;
assign a380 = ~a378 & ~a376;
assign a382 = ~i20 & i18;
assign a384 = a382 & i16;
assign a386 = a384 & ~i32;
assign a388 = ~a384 & i32;
assign a390 = ~a388 & ~a386;
assign a392 = ~i20 & ~i18;
assign a394 = a392 & ~i16;
assign a396 = a394 & ~i30;
assign a398 = ~a394 & i30;
assign a400 = ~a398 & ~a396;
assign a402 = a382 & ~i16;
assign a404 = a402 & ~i28;
assign a406 = ~a402 & i28;
assign a408 = ~a406 & ~a404;
assign a410 = a392 & i16;
assign a412 = a410 & ~i26;
assign a414 = ~a410 & i26;
assign a416 = ~a414 & ~a412;
assign a418 = i20 & ~i18;
assign a420 = a418 & i16;
assign a422 = ~a420 & i12;
assign a424 = a422 & ~i14;
assign a426 = ~a422 & i14;
assign a428 = ~a426 & ~a424;
assign a430 = ~i110 & ~i108;
assign a432 = a430 & ~i106;
assign a434 = a432 & ~i66;
assign a436 = i110 & i108;
assign a438 = a436 & ~i106;
assign a440 = a432 & i66;
assign a442 = ~i110 & i108;
assign a444 = a442 & ~i106;
assign a446 = i110 & ~i108;
assign a448 = a446 & i106;
assign a450 = ~a448 & ~a444;
assign a452 = a450 & ~a440;
assign a454 = a452 & ~a438;
assign a456 = ~a454 & i118;
assign a458 = ~a456 & ~a434;
assign a460 = ~a458 & ~i98;
assign a462 = a458 & i98;
assign a464 = ~a462 & ~a460;
assign a466 = a446 & ~i106;
assign a468 = a466 & i118;
assign a470 = a468 & ~a438;
assign a472 = ~a470 & i118;
assign a474 = a472 & a452;
assign a476 = ~a474 & ~a434;
assign a478 = a476 & ~i104;
assign a480 = ~a476 & i104;
assign a482 = ~a480 & ~a478;
assign a484 = ~a434 & ~i102;
assign a486 = a434 & i102;
assign a488 = ~a486 & ~a484;
assign a490 = a488 & a482;
assign a492 = i110 & ~i106;
assign a494 = ~a492 & a452;
assign a496 = ~a494 & i118;
assign a498 = ~a496 & ~a434;
assign a500 = a498 & ~i100;
assign a502 = ~a498 & i100;
assign a504 = ~a502 & ~a500;
assign a506 = a504 & a490;
assign a508 = ~a434 & ~i118;
assign a510 = a508 & ~i100;
assign a512 = ~a508 & i100;
assign a514 = ~a512 & ~a510;
assign a516 = ~a452 & i118;
assign a518 = ~a466 & i118;
assign a520 = a518 & ~a438;
assign a522 = a520 & ~a516;
assign a524 = ~a522 & ~a434;
assign a526 = a524 & ~i102;
assign a528 = ~a524 & i102;
assign a530 = ~a528 & ~a526;
assign a532 = a430 & ~i66;
assign a534 = a436 & i118;
assign a536 = a534 & a452;
assign a538 = ~a536 & ~a532;
assign a540 = ~a538 & ~i106;
assign a542 = ~a540 & ~i104;
assign a544 = a540 & i104;
assign a546 = ~a544 & ~a542;
assign a548 = a546 & a530;
assign a550 = ~a530 & ~a488;
assign a552 = ~a550 & a482;
assign a554 = ~a552 & ~a548;
assign a556 = ~a554 & a514;
assign a558 = ~a556 & ~a506;
assign a560 = ~a558 & ~i96;
assign a562 = a530 & a482;
assign a564 = a562 & a514;
assign a566 = a522 & ~a434;
assign a568 = a566 & ~i96;
assign a570 = ~a566 & i96;
assign a572 = ~a570 & ~a568;
assign a574 = a572 & a564;
assign a576 = ~a574 & ~a560;
assign a578 = ~a576 & a464;
assign a580 = a546 & a488;
assign a582 = a580 & a514;
assign a584 = a470 & a452;
assign a586 = ~a584 & i118;
assign a588 = ~a586 & ~a434;
assign a590 = ~a588 & ~i98;
assign a592 = a588 & i98;
assign a594 = ~a592 & ~a590;
assign a596 = a594 & a582;
assign a598 = a596 & ~i96;
assign a600 = a594 & a490;
assign a602 = a600 & a514;
assign a604 = a602 & ~i96;
assign a606 = a582 & a464;
assign a608 = a606 & ~i96;
assign a610 = a580 & a504;
assign a612 = a610 & a464;
assign a614 = a612 & ~i96;
assign a616 = a562 & a504;
assign a618 = a616 & a594;
assign a620 = a618 & ~i96;
assign a622 = a548 & a504;
assign a624 = a622 & a594;
assign a626 = a624 & ~i96;
assign a628 = a548 & a514;
assign a630 = a628 & a594;
assign a632 = a630 & ~i96;
assign a634 = a610 & a594;
assign a636 = a634 & ~i96;
assign a638 = a594 & a564;
assign a640 = a638 & ~i96;
assign a642 = a594 & a506;
assign a644 = a642 & ~i96;
assign a646 = a628 & a572;
assign a648 = a646 & a464;
assign a650 = a622 & a464;
assign a652 = a650 & ~i96;
assign a654 = a616 & a464;
assign a656 = a654 & ~i96;
assign a658 = ~a656 & ~a652;
assign a660 = a658 & ~a648;
assign a662 = a660 & ~a644;
assign a664 = a662 & ~a640;
assign a666 = a664 & ~a636;
assign a668 = a666 & ~a632;
assign a670 = a668 & ~a626;
assign a672 = a670 & ~a620;
assign a674 = a672 & ~a614;
assign a676 = a674 & ~a608;
assign a678 = a676 & ~a604;
assign a680 = a678 & ~a598;
assign a682 = a680 & ~a578;
assign a684 = ~a436 & ~i106;
assign a686 = ~a684 & ~a448;
assign a688 = a686 & ~a438;
assign a690 = ~i40 & ~i38;
assign a692 = i40 & i38;
assign a694 = ~a692 & ~a690;
assign a696 = ~a694 & i38;
assign a698 = ~a694 & i40;
assign a700 = i18 & ~i12;
assign a702 = ~i18 & i12;
assign a704 = ~a702 & ~a700;
assign a706 = i20 & ~i12;
assign a708 = ~i20 & i12;
assign a710 = ~a708 & ~a706;
assign a712 = a710 & a704;
assign a714 = ~a704 & i18;
assign a716 = ~a714 & ~i20;
assign a718 = ~a716 & ~a712;
assign a720 = ~a718 & ~i16;
assign a722 = i16 & ~i12;
assign a724 = ~i16 & i12;
assign a726 = ~a724 & ~a722;
assign a728 = a726 & a392;
assign a730 = a710 & ~i18;
assign a732 = a730 & a726;
assign a734 = a730 & ~i16;
assign a736 = a726 & a704;
assign a738 = a736 & ~i20;
assign a740 = ~a738 & ~a734;
assign a742 = a740 & ~a732;
assign a744 = a742 & ~a728;
assign a746 = a744 & ~a720;
assign a748 = ~a746 & ~a698;
assign a750 = a748 & ~a696;
assign a752 = a750 & ~a688;
assign a754 = a752 & ~a682;
assign a756 = a754 & i2;
assign a758 = a756 & ~i4;
assign a760 = a758 & i6;
assign a762 = a760 & ~i8;
assign a764 = a762 & ~i10;
assign a766 = a764 & a428;
assign a768 = ~a410 & ~a384;
assign a770 = a768 & ~a402;
assign a772 = a770 & ~a394;
assign a774 = ~a772 & ~i22;
assign a776 = a772 & i22;
assign a778 = ~a776 & ~a774;
assign a780 = a778 & a766;
assign a782 = a772 & ~a374;
assign a784 = a782 & a422;
assign a786 = a784 & ~i24;
assign a788 = ~a784 & i24;
assign a790 = ~a788 & ~a786;
assign a792 = a790 & a780;
assign a794 = a792 & a416;
assign a796 = a794 & a408;
assign a798 = a796 & a400;
assign a800 = a798 & a390;
assign a802 = a800 & a380;
assign a804 = a802 & ~i44;
assign a806 = a804 & ~i46;
assign a808 = a806 & a370;
assign a810 = a808 & i76;
assign a812 = a810 & i78;
assign a814 = a812 & ~i80;
assign a816 = a814 & ~i120;
assign a818 = a816 & ~i122;
assign a820 = a818 & i138;
assign a822 = a820 & ~i140;
assign a824 = a822 & ~i142;
assign a826 = a824 & ~i146;
assign a828 = a826 & ~i150;
assign a830 = a828 & ~i152;
assign a832 = a830 & ~i154;
assign a834 = a832 & ~i156;
assign a836 = a834 & ~i158;
assign a838 = a836 & ~i160;
assign a840 = a838 & ~i162;
assign a842 = ~a840 & ~l340;
assign a844 = ~l276 & ~l274;
assign a846 = a844 & ~l272;
assign a848 = a846 & ~l270;
assign a850 = a848 & ~l268;
assign a852 = a850 & ~l284;
assign a854 = a852 & i112;
assign a856 = a854 & l236;
assign a858 = a856 & ~l292;
assign a860 = a858 & l302;
assign a862 = ~l282 & l280;
assign a864 = a862 & ~l278;
assign a866 = a852 & l236;
assign a868 = a866 & ~a864;
assign a870 = a868 & ~l292;
assign a872 = a870 & l302;
assign a874 = a872 & ~l306;
assign a876 = a874 & i134;
assign a878 = a850 & l236;
assign a880 = a878 & ~l294;
assign a882 = a880 & l292;
assign a884 = a882 & l304;
assign a886 = a884 & ~l306;
assign a888 = a886 & i134;
assign a890 = a880 & ~a864;
assign a892 = a890 & a444;
assign a894 = a892 & l304;
assign a896 = a894 & l326;
assign a898 = a878 & ~i64;
assign a900 = a898 & ~l294;
assign a902 = a900 & l326;
assign a904 = a880 & l302;
assign a906 = a904 & ~i130;
assign a908 = a906 & l326;
assign a910 = a892 & ~l304;
assign a912 = a910 & l326;
assign a914 = a878 & ~a864;
assign a916 = a914 & ~i106;
assign a918 = a916 & ~i110;
assign a920 = a918 & i108;
assign a922 = a920 & l304;
assign a924 = a922 & l308;
assign a926 = a924 & ~l326;
assign a928 = a898 & ~l326;
assign a930 = a878 & l302;
assign a932 = a930 & ~i130;
assign a934 = a932 & ~l326;
assign a936 = a914 & ~i110;
assign a938 = a936 & i108;
assign a940 = a938 & ~i106;
assign a942 = a940 & ~l304;
assign a944 = a942 & ~l326;
assign a946 = a940 & ~l308;
assign a948 = a946 & ~l326;
assign a950 = l282 & l280;
assign a952 = a950 & ~l278;
assign a954 = ~a952 & a878;
assign a956 = a954 & a438;
assign a958 = l282 & ~l280;
assign a960 = a958 & ~l278;
assign a962 = ~a960 & a878;
assign a964 = a962 & a466;
assign a966 = a878 & l300;
assign a968 = a966 & ~i128;
assign a970 = a878 & l294;
assign a972 = a970 & ~a864;
assign a974 = a972 & ~i110;
assign a976 = a974 & i108;
assign a978 = a976 & ~i106;
assign a980 = a978 & l304;
assign a982 = a980 & l326;
assign a984 = a898 & l294;
assign a986 = a984 & l326;
assign a988 = a970 & l302;
assign a990 = a988 & ~i130;
assign a992 = a990 & l326;
assign a994 = a978 & ~l304;
assign a996 = a994 & l326;
assign a998 = ~l276 & l274;
assign a1000 = a998 & ~l272;
assign a1002 = a1000 & ~l270;
assign a1004 = a1002 & ~l268;
assign a1006 = a1004 & ~l284;
assign a1008 = a1006 & i112;
assign a1010 = a1008 & l236;
assign a1012 = a1004 & l236;
assign a1014 = a1012 & ~a864;
assign a1016 = a1014 & ~i110;
assign a1018 = a1016 & i108;
assign a1020 = a1018 & ~i106;
assign a1022 = a1020 & l302;
assign a1024 = a1022 & l304;
assign a1026 = a1006 & l236;
assign a1028 = a1026 & ~l292;
assign a1030 = a1028 & i120;
assign a1032 = a1012 & ~i64;
assign a1034 = a1012 & ~l292;
assign a1036 = a1034 & l302;
assign a1038 = a1036 & ~i130;
assign a1040 = a1020 & ~l304;
assign a1042 = a1012 & ~a952;
assign a1044 = a1042 & i110;
assign a1046 = a1044 & i108;
assign a1048 = a1046 & ~i106;
assign a1050 = a1012 & ~a960;
assign a1052 = a1050 & i110;
assign a1054 = a1052 & ~i108;
assign a1056 = a1054 & ~i106;
assign a1058 = a1012 & l300;
assign a1060 = a1058 & ~i128;
assign a1062 = a958 & l278;
assign a1064 = l276 & ~l274;
assign a1066 = a1064 & ~l272;
assign a1068 = a1066 & ~l270;
assign a1070 = a1068 & ~l268;
assign a1072 = a1070 & l236;
assign a1074 = a1072 & ~l294;
assign a1076 = a1074 & ~a1062;
assign a1078 = a1076 & a448;
assign a1080 = a1078 & ~l324;
assign a1082 = ~l282 & ~l280;
assign a1084 = a1082 & ~l278;
assign a1086 = ~a1084 & a1074;
assign a1088 = a1086 & a432;
assign a1090 = a1088 & ~l324;
assign a1092 = a1070 & ~l284;
assign a1094 = a1092 & i112;
assign a1096 = a1094 & l236;
assign a1098 = a1096 & a1062;
assign a1100 = a1098 & l302;
assign a1102 = a1096 & a1084;
assign a1104 = a1102 & l302;
assign a1106 = a1072 & ~a1062;
assign a1108 = a1106 & i110;
assign a1110 = a1108 & ~i108;
assign a1112 = a1110 & i106;
assign a1114 = a1112 & ~l292;
assign a1116 = a1114 & l324;
assign a1118 = ~a1084 & a1072;
assign a1120 = a1118 & ~i110;
assign a1122 = a1120 & ~i108;
assign a1124 = a1122 & ~i106;
assign a1126 = a1124 & ~l292;
assign a1128 = a1126 & l324;
assign a1130 = a1092 & l236;
assign a1132 = a1130 & a1062;
assign a1134 = a1132 & l292;
assign a1136 = a1134 & ~i120;
assign a1138 = a1136 & l302;
assign a1140 = a1138 & l324;
assign a1142 = a1130 & a1084;
assign a1144 = a1142 & l292;
assign a1146 = a1144 & ~i120;
assign a1148 = a1146 & l302;
assign a1150 = a1148 & l324;
assign a1152 = a1072 & ~i64;
assign a1154 = a1072 & l302;
assign a1156 = a1154 & ~i130;
assign a1158 = a1072 & a864;
assign a1160 = a1158 & l304;
assign a1162 = a1160 & ~i132;
assign a1164 = a1072 & ~a864;
assign a1166 = a1164 & ~i110;
assign a1168 = a1166 & i108;
assign a1170 = a1168 & ~i106;
assign a1172 = a1170 & ~l304;
assign a1174 = a1096 & a864;
assign a1176 = a1174 & l308;
assign a1178 = a1174 & ~l308;
assign a1180 = a1072 & ~a952;
assign a1182 = a1180 & i110;
assign a1184 = a1182 & i108;
assign a1186 = a1184 & ~i106;
assign a1188 = a1072 & ~a960;
assign a1190 = a1188 & i110;
assign a1192 = a1190 & ~i108;
assign a1194 = a1192 & ~i106;
assign a1196 = a1072 & l300;
assign a1198 = a1196 & ~i128;
assign a1200 = a1074 & i122;
assign a1202 = a998 & l272;
assign a1204 = a1202 & ~l270;
assign a1206 = a1204 & ~l268;
assign a1208 = a1206 & l236;
assign a1210 = a1208 & ~i64;
assign a1212 = a1210 & ~l238;
assign a1214 = a1212 & a1084;
assign a1216 = a1208 & a1084;
assign a1218 = a1216 & ~l302;
assign a1220 = a1218 & i130;
assign a1222 = a1220 & ~l324;
assign a1224 = a1208 & a1062;
assign a1226 = a1224 & ~l302;
assign a1228 = a1226 & i130;
assign a1230 = a1228 & ~l324;
assign a1232 = a1208 & ~a1084;
assign a1234 = a1232 & ~i110;
assign a1236 = a1234 & ~i108;
assign a1238 = a1236 & ~i106;
assign a1240 = a1238 & l302;
assign a1242 = a1240 & ~l324;
assign a1244 = a1208 & ~a1062;
assign a1246 = a1244 & i110;
assign a1248 = a1246 & ~i108;
assign a1250 = a1248 & i106;
assign a1252 = a1250 & l302;
assign a1254 = a1252 & ~l324;
assign a1256 = a1206 & ~l284;
assign a1258 = a1256 & l236;
assign a1260 = a1258 & a1084;
assign a1262 = a1260 & ~l292;
assign a1264 = a1262 & ~l302;
assign a1266 = a1264 & i130;
assign a1268 = a1266 & l324;
assign a1270 = a1258 & a1062;
assign a1272 = a1270 & ~l292;
assign a1274 = a1272 & ~l302;
assign a1276 = a1274 & i130;
assign a1278 = a1276 & l324;
assign a1280 = a1238 & ~l292;
assign a1282 = a1280 & l302;
assign a1284 = a1282 & l324;
assign a1286 = a1250 & ~l292;
assign a1288 = a1286 & l302;
assign a1290 = a1288 & l324;
assign a1292 = a1208 & ~l294;
assign a1294 = a1292 & ~a1084;
assign a1296 = a1294 & ~i110;
assign a1298 = a1296 & ~i108;
assign a1300 = a1298 & ~i106;
assign a1302 = a1300 & l292;
assign a1304 = a1302 & l302;
assign a1306 = a1304 & l324;
assign a1308 = a1292 & ~a1062;
assign a1310 = a1308 & i110;
assign a1312 = a1310 & ~i108;
assign a1314 = a1312 & i106;
assign a1316 = a1314 & l292;
assign a1318 = a1316 & l302;
assign a1320 = a1318 & l324;
assign a1322 = a1258 & ~l294;
assign a1324 = a1322 & a1084;
assign a1326 = a1324 & l292;
assign a1328 = a1326 & ~l302;
assign a1330 = a1328 & i130;
assign a1332 = a1322 & a1062;
assign a1334 = a1332 & l292;
assign a1336 = a1334 & ~l302;
assign a1338 = a1336 & i130;
assign a1340 = a1322 & a864;
assign a1342 = a1340 & ~l302;
assign a1344 = a1342 & i130;
assign a1346 = a1344 & l304;
assign a1348 = a1340 & l302;
assign a1350 = a1348 & ~l304;
assign a1352 = a1350 & i132;
assign a1354 = a1256 & i112;
assign a1356 = a1354 & l236;
assign a1358 = a1208 & ~a952;
assign a1360 = a1358 & i110;
assign a1362 = a1360 & i108;
assign a1364 = a1362 & ~i106;
assign a1366 = a1208 & ~a960;
assign a1368 = a1366 & i110;
assign a1370 = a1368 & ~i108;
assign a1372 = a1370 & ~i106;
assign a1374 = a1208 & l300;
assign a1376 = a1374 & ~i128;
assign a1378 = a1292 & i122;
assign a1380 = a1206 & ~l236;
assign a1382 = a1380 & ~l238;
assign a1384 = a1382 & ~a1084;
assign a1386 = a1384 & ~i110;
assign a1388 = a1386 & ~i108;
assign a1390 = a1388 & ~i106;
assign a1392 = a1390 & ~l314;
assign a1394 = a1354 & ~l236;
assign a1396 = a1394 & ~l238;
assign a1398 = a1396 & a1084;
assign a1400 = a1394 & l238;
assign a1402 = a1400 & a1084;
assign a1404 = a1402 & l296;
assign a1406 = a1390 & l314;
assign a1408 = a1406 & ~l310;
assign a1410 = a1380 & ~l216;
assign a1412 = a1410 & i44;
assign a1414 = a1412 & ~l238;
assign a1416 = a1394 & a1062;
assign a1418 = a1394 & a864;
assign a1420 = a1402 & ~l296;
assign a1422 = a1380 & ~a952;
assign a1424 = a1422 & i110;
assign a1426 = a1424 & i108;
assign a1428 = a1426 & ~i106;
assign a1430 = a1380 & ~a960;
assign a1432 = a1430 & i110;
assign a1434 = a1432 & ~i108;
assign a1436 = a1434 & ~i106;
assign a1438 = a1380 & ~l288;
assign a1440 = a1438 & l290;
assign a1442 = a1440 & ~i118;
assign a1444 = a1380 & ~l294;
assign a1446 = a1444 & i122;
assign a1448 = a1438 & i116;
assign a1450 = a848 & l268;
assign a1452 = a1450 & l236;
assign a1454 = a1452 & ~a1062;
assign a1456 = a1454 & i110;
assign a1458 = a1456 & ~i108;
assign a1460 = a1458 & i106;
assign a1462 = a1460 & l302;
assign a1464 = a1452 & ~a1084;
assign a1466 = a1464 & ~i110;
assign a1468 = a1466 & ~i108;
assign a1470 = a1468 & ~i106;
assign a1472 = a1470 & l302;
assign a1474 = a1464 & l308;
assign a1476 = a1474 & ~i136;
assign a1478 = a1452 & ~i64;
assign a1480 = a1452 & l302;
assign a1482 = a1480 & ~i130;
assign a1484 = a1452 & l304;
assign a1486 = a1484 & ~i132;
assign a1488 = a1452 & ~a952;
assign a1490 = a1488 & i110;
assign a1492 = a1490 & i108;
assign a1494 = a1492 & ~i106;
assign a1496 = a1452 & ~a960;
assign a1498 = a1496 & i110;
assign a1500 = a1498 & ~i108;
assign a1502 = a1500 & ~i106;
assign a1504 = a1452 & l300;
assign a1506 = a1504 & ~i128;
assign a1508 = l276 & l274;
assign a1510 = a1508 & ~l272;
assign a1512 = a1510 & l270;
assign a1514 = a1512 & ~l268;
assign a1516 = a1514 & l236;
assign a1518 = a1516 & a1084;
assign a1520 = a1518 & ~l302;
assign a1522 = a1520 & i130;
assign a1524 = a1516 & a1062;
assign a1526 = a1524 & ~l302;
assign a1528 = a1526 & i130;
assign a1530 = a1516 & ~a1084;
assign a1532 = a1530 & ~i110;
assign a1534 = a1532 & ~i108;
assign a1536 = a1534 & ~i106;
assign a1538 = a1536 & l302;
assign a1540 = a1516 & ~a1062;
assign a1542 = a1540 & i110;
assign a1544 = a1542 & ~i108;
assign a1546 = a1544 & i106;
assign a1548 = a1546 & l302;
assign a1550 = a1516 & a864;
assign a1552 = a1550 & ~l302;
assign a1554 = a1552 & i130;
assign a1556 = a1554 & l304;
assign a1558 = a1556 & l308;
assign a1560 = a1550 & l302;
assign a1562 = a1560 & ~l304;
assign a1564 = a1562 & i132;
assign a1566 = a1564 & l308;
assign a1568 = a1516 & l302;
assign a1570 = a1568 & l304;
assign a1572 = a1570 & ~l308;
assign a1574 = a1572 & i136;
assign a1576 = a1516 & ~a952;
assign a1578 = a1576 & i110;
assign a1580 = a1578 & i108;
assign a1582 = a1580 & ~i106;
assign a1584 = a1516 & ~a960;
assign a1586 = a1584 & i110;
assign a1588 = a1586 & ~i108;
assign a1590 = a1588 & ~i106;
assign a1592 = a1516 & l300;
assign a1594 = a1592 & ~i128;
assign a1596 = a1514 & ~l236;
assign a1598 = a1596 & ~l238;
assign a1600 = a1598 & ~a1084;
assign a1602 = a1600 & ~i110;
assign a1604 = a1602 & ~i108;
assign a1606 = a1604 & ~i106;
assign a1608 = a1514 & ~l284;
assign a1610 = a1608 & i112;
assign a1612 = a1610 & ~l236;
assign a1614 = a1612 & l238;
assign a1616 = a1614 & a1084;
assign a1618 = a1616 & l296;
assign a1620 = a1596 & ~l216;
assign a1622 = a1620 & i44;
assign a1624 = a1622 & ~l238;
assign a1626 = a1596 & ~a952;
assign a1628 = a1626 & i110;
assign a1630 = a1628 & i108;
assign a1632 = a1630 & ~i106;
assign a1634 = a1596 & ~a960;
assign a1636 = a1634 & i110;
assign a1638 = a1636 & ~i108;
assign a1640 = a1638 & ~i106;
assign a1642 = a1596 & ~l288;
assign a1644 = a1642 & l290;
assign a1646 = a1644 & ~i118;
assign a1648 = a1642 & i116;
assign a1650 = a1000 & l270;
assign a1652 = a1650 & ~l268;
assign a1654 = a1652 & l236;
assign a1656 = a1654 & ~a1084;
assign a1658 = a1656 & ~i110;
assign a1660 = a1658 & ~i108;
assign a1662 = a1660 & ~i106;
assign a1664 = a1662 & l302;
assign a1666 = a1654 & ~a1062;
assign a1668 = a1666 & i110;
assign a1670 = a1668 & ~i108;
assign a1672 = a1670 & i106;
assign a1674 = a1672 & l302;
assign a1676 = a1654 & ~a864;
assign a1678 = a1676 & ~i106;
assign a1680 = a1678 & ~i110;
assign a1682 = a1680 & i108;
assign a1684 = a1682 & l302;
assign a1686 = a1684 & l304;
assign a1688 = a1686 & l308;
assign a1690 = a1676 & ~i110;
assign a1692 = a1690 & i108;
assign a1694 = a1692 & ~i106;
assign a1696 = a1694 & ~l302;
assign a1698 = a1694 & ~l304;
assign a1700 = a1694 & ~l308;
assign a1702 = a1662 & ~l302;
assign a1704 = a1672 & ~l302;
assign a1706 = a1654 & ~a960;
assign a1708 = a1706 & i110;
assign a1710 = a1708 & ~i108;
assign a1712 = a1710 & ~i106;
assign a1714 = a1654 & l300;
assign a1716 = a1714 & ~i128;
assign a1718 = a1652 & ~l236;
assign a1720 = a1718 & ~l238;
assign a1722 = a1720 & ~a1084;
assign a1724 = a1722 & ~i110;
assign a1726 = a1724 & ~i108;
assign a1728 = a1726 & ~i106;
assign a1730 = a1718 & ~a864;
assign a1732 = a1730 & ~i110;
assign a1734 = a1732 & i108;
assign a1736 = a1734 & ~i106;
assign a1738 = a1718 & ~a1062;
assign a1740 = a1738 & i110;
assign a1742 = a1740 & ~i108;
assign a1744 = a1742 & i106;
assign a1746 = a1718 & l238;
assign a1748 = a1746 & ~a1084;
assign a1750 = a1748 & ~i110;
assign a1752 = a1750 & ~i108;
assign a1754 = a1752 & ~i106;
assign a1756 = a1718 & ~a960;
assign a1758 = a1756 & i110;
assign a1760 = a1758 & ~i108;
assign a1762 = a1760 & ~i106;
assign a1764 = a1718 & ~l288;
assign a1766 = a1764 & l290;
assign a1768 = a1766 & ~i118;
assign a1770 = a1764 & i116;
assign a1772 = a1510 & ~l270;
assign a1774 = a1772 & ~l268;
assign a1776 = a1774 & l236;
assign a1778 = a1776 & ~a1084;
assign a1780 = a1778 & ~i110;
assign a1782 = a1780 & ~i108;
assign a1784 = a1782 & ~i106;
assign a1786 = a1784 & l302;
assign a1788 = a1776 & ~a1062;
assign a1790 = a1788 & i110;
assign a1792 = a1790 & ~i108;
assign a1794 = a1792 & i106;
assign a1796 = a1794 & l302;
assign a1798 = a1776 & ~a864;
assign a1800 = a1798 & ~i106;
assign a1802 = a1800 & ~i110;
assign a1804 = a1802 & i108;
assign a1806 = a1804 & l302;
assign a1808 = a1806 & l304;
assign a1810 = a1808 & l308;
assign a1812 = a1798 & ~i110;
assign a1814 = a1812 & i108;
assign a1816 = a1814 & ~i106;
assign a1818 = a1816 & ~l302;
assign a1820 = a1816 & ~l304;
assign a1822 = a1816 & ~l308;
assign a1824 = a1784 & ~l302;
assign a1826 = a1794 & ~l302;
assign a1828 = a1776 & ~a952;
assign a1830 = a1828 & i110;
assign a1832 = a1830 & i108;
assign a1834 = a1832 & ~i106;
assign a1836 = a1776 & l300;
assign a1838 = a1836 & ~i128;
assign a1840 = a1774 & ~l236;
assign a1842 = a1840 & ~l238;
assign a1844 = a1842 & ~a1084;
assign a1846 = a1844 & ~i110;
assign a1848 = a1846 & ~i108;
assign a1850 = a1848 & ~i106;
assign a1852 = a1840 & ~a864;
assign a1854 = a1852 & ~i110;
assign a1856 = a1854 & i108;
assign a1858 = a1856 & ~i106;
assign a1860 = a1840 & ~a1062;
assign a1862 = a1860 & i110;
assign a1864 = a1862 & ~i108;
assign a1866 = a1864 & i106;
assign a1868 = a1840 & l238;
assign a1870 = a1868 & ~a1084;
assign a1872 = a1870 & ~i110;
assign a1874 = a1872 & ~i108;
assign a1876 = a1874 & ~i106;
assign a1878 = a1840 & ~a952;
assign a1880 = a1878 & i110;
assign a1882 = a1880 & i108;
assign a1884 = a1882 & ~i106;
assign a1886 = a1840 & ~l288;
assign a1888 = a1886 & l290;
assign a1890 = a1888 & ~i118;
assign a1892 = a1886 & i116;
assign a1894 = a1508 & l272;
assign a1896 = a1894 & ~l270;
assign a1898 = a1896 & ~l268;
assign a1900 = a1898 & l236;
assign a1902 = a1900 & a1084;
assign a1904 = a1902 & ~l300;
assign a1906 = a1904 & i128;
assign a1908 = a1906 & l302;
assign a1910 = a1900 & a1062;
assign a1912 = a1910 & ~l300;
assign a1914 = a1912 & i128;
assign a1916 = a1914 & l302;
assign a1918 = a1900 & a864;
assign a1920 = a1918 & ~l300;
assign a1922 = a1920 & i128;
assign a1924 = a1922 & l302;
assign a1926 = a1924 & l304;
assign a1928 = a1926 & l308;
assign a1930 = a1922 & ~l302;
assign a1932 = a1922 & ~l304;
assign a1934 = a1922 & ~l308;
assign a1936 = a1906 & ~l302;
assign a1938 = a1914 & ~l302;
assign a1940 = a1900 & a952;
assign a1942 = a1940 & ~l300;
assign a1944 = a1942 & i128;
assign a1946 = a1900 & a960;
assign a1948 = a1946 & ~l300;
assign a1950 = a1948 & i128;
assign a1952 = a1898 & ~l236;
assign a1954 = a1952 & ~l238;
assign a1956 = a1954 & ~l290;
assign a1958 = a1956 & i118;
assign a1960 = a1958 & a1084;
assign a1962 = a1952 & ~l290;
assign a1964 = a1962 & i118;
assign a1966 = a1964 & a864;
assign a1968 = a1964 & a1062;
assign a1970 = a1952 & l238;
assign a1972 = a1970 & ~l290;
assign a1974 = a1972 & i118;
assign a1976 = a1974 & a1084;
assign a1978 = a1964 & a952;
assign a1980 = a1964 & a960;
assign a1982 = a1952 & ~l288;
assign a1984 = a1982 & i116;
assign a1986 = a844 & l272;
assign a1988 = a1986 & l270;
assign a1990 = a1988 & ~l268;
assign a1992 = a1990 & ~l284;
assign a1994 = a1992 & i112;
assign a1996 = a1994 & l236;
assign a1998 = a1996 & a1062;
assign a2000 = a1998 & l302;
assign a2002 = a1996 & a1084;
assign a2004 = a2002 & l302;
assign a2006 = a1996 & a864;
assign a2008 = a2006 & l308;
assign a2010 = a2006 & ~l308;
assign a2012 = a1990 & l236;
assign a2014 = a2012 & ~a952;
assign a2016 = a2014 & i110;
assign a2018 = a2016 & i108;
assign a2020 = a2018 & ~i106;
assign a2022 = a2012 & ~a960;
assign a2024 = a2022 & i110;
assign a2026 = a2024 & ~i108;
assign a2028 = a2026 & ~i106;
assign a2030 = a2012 & l300;
assign a2032 = a2030 & ~i128;
assign a2034 = a2012 & l302;
assign a2036 = a2034 & ~i130;
assign a2038 = a2012 & a864;
assign a2040 = a2038 & l304;
assign a2042 = a2040 & ~i132;
assign a2044 = a2012 & ~a864;
assign a2046 = a2044 & ~i110;
assign a2048 = a2046 & i108;
assign a2050 = a2048 & ~i106;
assign a2052 = a2050 & ~l304;
assign a2054 = a2012 & ~i64;
assign a2056 = a1064 & l272;
assign a2058 = a2056 & l270;
assign a2060 = a2058 & ~l268;
assign a2062 = a2060 & l236;
assign a2064 = a2062 & ~i64;
assign a2066 = a2064 & ~l238;
assign a2068 = a2066 & a1084;
assign a2070 = a2062 & a1084;
assign a2072 = a2070 & ~l302;
assign a2074 = a2072 & i130;
assign a2076 = a2074 & ~l324;
assign a2078 = a2062 & a1062;
assign a2080 = a2078 & ~l302;
assign a2082 = a2080 & i130;
assign a2084 = a2082 & ~l324;
assign a2086 = a2062 & ~a1084;
assign a2088 = a2086 & ~i110;
assign a2090 = a2088 & ~i108;
assign a2092 = a2090 & ~i106;
assign a2094 = a2092 & l302;
assign a2096 = a2094 & ~l324;
assign a2098 = a2062 & ~a1062;
assign a2100 = a2098 & i110;
assign a2102 = a2100 & ~i108;
assign a2104 = a2102 & i106;
assign a2106 = a2104 & l302;
assign a2108 = a2106 & ~l324;
assign a2110 = a2060 & ~l284;
assign a2112 = a2110 & i112;
assign a2114 = a2112 & l236;
assign a2116 = a2114 & a1084;
assign a2118 = a2116 & l302;
assign a2120 = a2114 & a1062;
assign a2122 = a2120 & l302;
assign a2124 = a2114 & a864;
assign a2126 = a2114 & ~l302;
assign a2128 = a2062 & ~a952;
assign a2130 = a2128 & i110;
assign a2132 = a2130 & i108;
assign a2134 = a2132 & ~i106;
assign a2136 = a2062 & ~a960;
assign a2138 = a2136 & i110;
assign a2140 = a2138 & ~i108;
assign a2142 = a2140 & ~i106;
assign a2144 = a2062 & l300;
assign a2146 = a2144 & ~i128;
assign a2148 = a2062 & a864;
assign a2150 = a2148 & ~l302;
assign a2152 = a2150 & i130;
assign a2154 = a2152 & l304;
assign a2156 = a2074 & l324;
assign a2158 = a2082 & l324;
assign a2160 = a2078 & l302;
assign a2162 = a2160 & ~l304;
assign a2164 = a2162 & i132;
assign a2166 = a2094 & l324;
assign a2168 = a2106 & l324;
assign a2170 = a2060 & ~l236;
assign a2172 = a2170 & ~l238;
assign a2174 = a2172 & ~a1084;
assign a2176 = a2174 & ~i110;
assign a2178 = a2176 & ~i108;
assign a2180 = a2178 & ~i106;
assign a2182 = a2180 & l310;
assign a2184 = a2112 & ~l236;
assign a2186 = a2184 & ~l238;
assign a2188 = a2186 & a1084;
assign a2190 = a2184 & l238;
assign a2192 = a2190 & a1084;
assign a2194 = a2192 & l296;
assign a2196 = a2180 & l314;
assign a2198 = a2196 & ~l310;
assign a2200 = a2170 & ~l216;
assign a2202 = a2200 & i44;
assign a2204 = a2202 & ~l238;
assign a2206 = a2184 & a1062;
assign a2208 = a2184 & a864;
assign a2210 = a2192 & ~l296;
assign a2212 = a2170 & ~a952;
assign a2214 = a2212 & i110;
assign a2216 = a2214 & i108;
assign a2218 = a2216 & ~i106;
assign a2220 = a2170 & ~a960;
assign a2222 = a2220 & i110;
assign a2224 = a2222 & ~i108;
assign a2226 = a2224 & ~i106;
assign a2228 = a2170 & ~l288;
assign a2230 = a2228 & l290;
assign a2232 = a2230 & ~i118;
assign a2234 = a2228 & i116;
assign a2236 = a1066 & l270;
assign a2238 = a2236 & ~l268;
assign a2240 = a2238 & ~l284;
assign a2242 = a2240 & i112;
assign a2244 = a2242 & ~l236;
assign a2246 = a2244 & a1084;
assign a2248 = a2238 & ~l236;
assign a2250 = a2248 & ~l288;
assign a2252 = a2250 & ~l294;
assign a2254 = a2252 & ~l328;
assign a2256 = a2254 & i154;
assign a2258 = a2248 & ~a1062;
assign a2260 = a2258 & i110;
assign a2262 = a2260 & ~i108;
assign a2264 = a2262 & i106;
assign a2266 = a2248 & ~a864;
assign a2268 = a2266 & ~i110;
assign a2270 = a2268 & i108;
assign a2272 = a2270 & ~i106;
assign a2274 = a2248 & i64;
assign a2276 = a2248 & ~a952;
assign a2278 = a2276 & i110;
assign a2280 = a2278 & i108;
assign a2282 = a2280 & ~i106;
assign a2284 = a2248 & ~a960;
assign a2286 = a2284 & i110;
assign a2288 = a2286 & ~i108;
assign a2290 = a2288 & ~i106;
assign a2292 = a2250 & l290;
assign a2294 = a2292 & ~i118;
assign a2296 = a2250 & l294;
assign a2298 = a2296 & ~l328;
assign a2300 = a2298 & i154;
assign a2302 = a2250 & i116;
assign a2304 = a1894 & l270;
assign a2306 = a2304 & ~l268;
assign a2308 = a2306 & ~l284;
assign a2310 = a2308 & i112;
assign a2312 = a2310 & ~l236;
assign a2314 = a2312 & a1084;
assign a2316 = a2306 & ~l236;
assign a2318 = a2316 & ~l288;
assign a2320 = a2318 & ~l294;
assign a2322 = a2320 & ~l328;
assign a2324 = a2322 & i154;
assign a2326 = a2316 & ~a1062;
assign a2328 = a2326 & i110;
assign a2330 = a2328 & ~i108;
assign a2332 = a2330 & i106;
assign a2334 = a2316 & ~a864;
assign a2336 = a2334 & ~i110;
assign a2338 = a2336 & i108;
assign a2340 = a2338 & ~i106;
assign a2342 = a2316 & i64;
assign a2344 = a2308 & ~l236;
assign a2346 = a2344 & ~l288;
assign a2348 = a2346 & l296;
assign a2350 = a2348 & ~i124;
assign a2352 = a2350 & ~l328;
assign a2354 = a2316 & ~a952;
assign a2356 = a2354 & i110;
assign a2358 = a2356 & i108;
assign a2360 = a2358 & ~i106;
assign a2362 = a2316 & ~a960;
assign a2364 = a2362 & i110;
assign a2366 = a2364 & ~i108;
assign a2368 = a2366 & ~i106;
assign a2370 = a2318 & l290;
assign a2372 = a2370 & ~i118;
assign a2374 = a2318 & l294;
assign a2376 = a2374 & ~l328;
assign a2378 = a2376 & i154;
assign a2380 = a2318 & i116;
assign a2382 = a846 & l270;
assign a2384 = a2382 & ~l268;
assign a2386 = a2384 & ~l236;
assign a2388 = a2386 & ~l286;
assign a2390 = a2388 & i114;
assign a2392 = a2390 & l314;
assign a2394 = a2384 & ~l284;
assign a2396 = a2394 & i112;
assign a2398 = a2396 & ~l236;
assign a2400 = a2386 & ~l216;
assign a2402 = a2400 & i44;
assign a2404 = a2386 & i64;
assign a2406 = a2404 & ~l294;
assign a2408 = a2406 & l326;
assign a2410 = a2386 & ~l238;
assign a2412 = a2410 & i66;
assign a2414 = a2412 & ~l294;
assign a2416 = a2414 & l326;
assign a2418 = a2386 & ~l294;
assign a2420 = a2418 & ~a864;
assign a2422 = a2420 & ~i110;
assign a2424 = a2422 & i108;
assign a2426 = a2424 & ~i106;
assign a2428 = a2426 & l326;
assign a2430 = a2418 & ~a1062;
assign a2432 = a2430 & i110;
assign a2434 = a2432 & ~i108;
assign a2436 = a2434 & i106;
assign a2438 = a2436 & l326;
assign a2440 = a2386 & ~a864;
assign a2442 = a2440 & ~i110;
assign a2444 = a2442 & i108;
assign a2446 = a2444 & ~i106;
assign a2448 = a2446 & ~l326;
assign a2450 = a2386 & ~a1062;
assign a2452 = a2450 & i110;
assign a2454 = a2452 & ~i108;
assign a2456 = a2454 & i106;
assign a2458 = a2456 & ~l326;
assign a2460 = a2412 & ~l326;
assign a2462 = a2404 & ~l326;
assign a2464 = a2386 & ~a952;
assign a2466 = a2464 & i110;
assign a2468 = a2466 & i108;
assign a2470 = a2468 & ~i106;
assign a2472 = a2386 & ~a960;
assign a2474 = a2472 & i110;
assign a2476 = a2474 & ~i108;
assign a2478 = a2476 & ~i106;
assign a2480 = a2386 & ~l288;
assign a2482 = a2480 & l290;
assign a2484 = a2482 & ~i118;
assign a2486 = a2404 & l294;
assign a2488 = a2486 & l326;
assign a2490 = a2412 & l294;
assign a2492 = a2490 & l326;
assign a2494 = a2386 & l294;
assign a2496 = a2494 & ~a864;
assign a2498 = a2496 & ~i110;
assign a2500 = a2498 & i108;
assign a2502 = a2500 & ~i106;
assign a2504 = a2502 & l326;
assign a2506 = a2494 & ~a1062;
assign a2508 = a2506 & i110;
assign a2510 = a2508 & ~i108;
assign a2512 = a2510 & i106;
assign a2514 = a2512 & l326;
assign a2516 = a2480 & i116;
assign a2518 = a1202 & l270;
assign a2520 = a2518 & ~l268;
assign a2522 = a2520 & ~l236;
assign a2524 = a2522 & ~l286;
assign a2526 = a2524 & i114;
assign a2528 = a2526 & l238;
assign a2530 = a2528 & ~l288;
assign a2532 = a2530 & l318;
assign a2534 = a2522 & l238;
assign a2536 = a2534 & ~i66;
assign a2538 = a2536 & ~l288;
assign a2540 = a2520 & ~l284;
assign a2542 = a2540 & i112;
assign a2544 = a2542 & ~l236;
assign a2546 = a2522 & i64;
assign a2548 = a2546 & ~l294;
assign a2550 = a2548 & l326;
assign a2552 = a2534 & ~l288;
assign a2554 = a2552 & ~l294;
assign a2556 = a2554 & ~a952;
assign a2558 = a2556 & ~a960;
assign a2560 = a2558 & l296;
assign a2562 = a2560 & ~i124;
assign a2564 = a2562 & l326;
assign a2566 = a2522 & ~l294;
assign a2568 = a2566 & ~a864;
assign a2570 = a2568 & ~i110;
assign a2572 = a2570 & i108;
assign a2574 = a2572 & ~i106;
assign a2576 = a2574 & l326;
assign a2578 = a2566 & ~a1062;
assign a2580 = a2578 & i110;
assign a2582 = a2580 & ~i108;
assign a2584 = a2582 & i106;
assign a2586 = a2584 & l326;
assign a2588 = a2522 & ~a864;
assign a2590 = a2588 & ~i110;
assign a2592 = a2590 & i108;
assign a2594 = a2592 & ~i106;
assign a2596 = a2594 & ~l326;
assign a2598 = a2522 & ~a1062;
assign a2600 = a2598 & i110;
assign a2602 = a2600 & ~i108;
assign a2604 = a2602 & i106;
assign a2606 = a2604 & ~l326;
assign a2608 = a2552 & ~a952;
assign a2610 = a2608 & ~a960;
assign a2612 = a2610 & l296;
assign a2614 = a2612 & ~i124;
assign a2616 = a2614 & ~l326;
assign a2618 = a2546 & ~l326;
assign a2620 = a2522 & ~a952;
assign a2622 = a2620 & i110;
assign a2624 = a2622 & i108;
assign a2626 = a2624 & ~i106;
assign a2628 = a2522 & ~a960;
assign a2630 = a2628 & i110;
assign a2632 = a2630 & ~i108;
assign a2634 = a2632 & ~i106;
assign a2636 = a2522 & ~l288;
assign a2638 = a2636 & l290;
assign a2640 = a2638 & ~i118;
assign a2642 = a2546 & l294;
assign a2644 = a2642 & l326;
assign a2646 = a2552 & l294;
assign a2648 = a2646 & ~a952;
assign a2650 = a2648 & ~a960;
assign a2652 = a2650 & l296;
assign a2654 = a2652 & ~i124;
assign a2656 = a2654 & l326;
assign a2658 = a2522 & l294;
assign a2660 = a2658 & ~a864;
assign a2662 = a2660 & ~i110;
assign a2664 = a2662 & i108;
assign a2666 = a2664 & ~i106;
assign a2668 = a2666 & l326;
assign a2670 = a2658 & ~a1062;
assign a2672 = a2670 & i110;
assign a2674 = a2672 & ~i108;
assign a2676 = a2674 & i106;
assign a2678 = a2676 & l326;
assign a2680 = a2636 & i116;
assign a2682 = a1068 & l268;
assign a2684 = a2682 & ~l236;
assign a2686 = a2684 & ~l286;
assign a2688 = a2686 & i114;
assign a2690 = a2682 & ~l284;
assign a2692 = a2690 & i112;
assign a2694 = a2692 & ~l236;
assign a2696 = a2684 & ~l216;
assign a2698 = a2696 & i44;
assign a2700 = a2684 & i64;
assign a2702 = a2700 & ~l294;
assign a2704 = a2684 & ~l294;
assign a2706 = a2704 & ~a864;
assign a2708 = a2706 & ~i110;
assign a2710 = a2708 & i108;
assign a2712 = a2710 & ~i106;
assign a2714 = a2704 & ~a1062;
assign a2716 = a2714 & i110;
assign a2718 = a2716 & ~i108;
assign a2720 = a2718 & i106;
assign a2722 = a2684 & ~a952;
assign a2724 = a2722 & i110;
assign a2726 = a2724 & i108;
assign a2728 = a2726 & ~i106;
assign a2730 = a2684 & ~a960;
assign a2732 = a2730 & i110;
assign a2734 = a2732 & ~i108;
assign a2736 = a2734 & ~i106;
assign a2738 = a2684 & ~l288;
assign a2740 = a2738 & l290;
assign a2742 = a2740 & ~i118;
assign a2744 = a2700 & l294;
assign a2746 = a2684 & l294;
assign a2748 = a2746 & ~a864;
assign a2750 = a2748 & ~i110;
assign a2752 = a2750 & i108;
assign a2754 = a2752 & ~i106;
assign a2756 = a2746 & ~a1062;
assign a2758 = a2756 & i110;
assign a2760 = a2758 & ~i108;
assign a2762 = a2760 & i106;
assign a2764 = a2738 & i116;
assign a2766 = ~a2764 & l268;
assign a2768 = a2766 & ~a2762;
assign a2770 = a2768 & ~a2754;
assign a2772 = a2770 & ~a2744;
assign a2774 = a2772 & ~a2742;
assign a2776 = a2774 & ~a2736;
assign a2778 = a2776 & ~a2728;
assign a2780 = a2778 & ~a2720;
assign a2782 = a2780 & ~a2712;
assign a2784 = a2782 & ~a2702;
assign a2786 = a2784 & ~a2698;
assign a2788 = a2786 & ~a2694;
assign a2790 = a2788 & ~a2688;
assign a2792 = a2790 & ~a2680;
assign a2794 = a2792 & ~a2678;
assign a2796 = a2794 & ~a2668;
assign a2798 = a2796 & ~a2656;
assign a2800 = a2798 & ~a2644;
assign a2802 = a2800 & ~a2640;
assign a2804 = a2802 & ~a2634;
assign a2806 = a2804 & ~a2626;
assign a2808 = a2806 & ~a2618;
assign a2810 = a2808 & ~a2616;
assign a2812 = a2810 & ~a2606;
assign a2814 = a2812 & ~a2596;
assign a2816 = a2814 & ~a2586;
assign a2818 = a2816 & ~a2576;
assign a2820 = a2818 & ~a2564;
assign a2822 = a2820 & ~a2550;
assign a2824 = a2822 & ~a2544;
assign a2826 = a2824 & ~a2538;
assign a2828 = a2826 & ~a2532;
assign a2830 = a2828 & ~a2516;
assign a2832 = a2830 & ~a2514;
assign a2834 = a2832 & ~a2504;
assign a2836 = a2834 & ~a2492;
assign a2838 = a2836 & ~a2488;
assign a2840 = a2838 & ~a2484;
assign a2842 = a2840 & ~a2478;
assign a2844 = a2842 & ~a2470;
assign a2846 = a2844 & ~a2462;
assign a2848 = a2846 & ~a2460;
assign a2850 = a2848 & ~a2458;
assign a2852 = a2850 & ~a2448;
assign a2854 = a2852 & ~a2438;
assign a2856 = a2854 & ~a2428;
assign a2858 = a2856 & ~a2416;
assign a2860 = a2858 & ~a2408;
assign a2862 = a2860 & ~a2402;
assign a2864 = a2862 & ~a2398;
assign a2866 = a2864 & ~a2392;
assign a2868 = a2866 & ~a2380;
assign a2870 = a2868 & ~a2378;
assign a2872 = a2870 & ~a2372;
assign a2874 = a2872 & ~a2368;
assign a2876 = a2874 & ~a2360;
assign a2878 = a2876 & ~a2352;
assign a2880 = a2878 & ~a2342;
assign a2882 = a2880 & ~a2340;
assign a2884 = a2882 & ~a2332;
assign a2886 = a2884 & ~a2324;
assign a2888 = a2886 & ~a2314;
assign a2890 = a2888 & ~a2302;
assign a2892 = a2890 & ~a2300;
assign a2894 = a2892 & ~a2294;
assign a2896 = a2894 & ~a2290;
assign a2898 = a2896 & ~a2282;
assign a2900 = a2898 & ~a2274;
assign a2902 = a2900 & ~a2272;
assign a2904 = a2902 & ~a2264;
assign a2906 = a2904 & ~a2256;
assign a2908 = a2906 & ~a2246;
assign a2910 = a2908 & ~a2234;
assign a2912 = a2910 & ~a2232;
assign a2914 = a2912 & ~a2226;
assign a2916 = a2914 & ~a2218;
assign a2918 = a2916 & ~a2210;
assign a2920 = a2918 & ~a2208;
assign a2922 = a2920 & ~a2206;
assign a2924 = a2922 & ~a2204;
assign a2926 = ~a2924 & ~a2198;
assign a2928 = ~a2926 & ~a2194;
assign a2930 = a2928 & ~a2188;
assign a2932 = a2930 & ~a2182;
assign a2934 = a2932 & ~a2168;
assign a2936 = a2934 & ~a2166;
assign a2938 = a2936 & ~a2164;
assign a2940 = a2938 & ~a2158;
assign a2942 = a2940 & ~a2156;
assign a2944 = a2942 & ~a2154;
assign a2946 = a2944 & ~a2146;
assign a2948 = a2946 & ~a2142;
assign a2950 = a2948 & ~a2134;
assign a2952 = a2950 & ~a2126;
assign a2954 = a2952 & ~a2124;
assign a2956 = a2954 & ~a2122;
assign a2958 = a2956 & ~a2118;
assign a2960 = a2958 & ~a2108;
assign a2962 = a2960 & ~a2096;
assign a2964 = a2962 & ~a2084;
assign a2966 = a2964 & ~a2076;
assign a2968 = a2966 & ~a2068;
assign a2970 = a2968 & ~a2054;
assign a2972 = a2970 & ~a2052;
assign a2974 = a2972 & ~a2042;
assign a2976 = a2974 & ~a2036;
assign a2978 = a2976 & ~a2032;
assign a2980 = a2978 & ~a2028;
assign a2982 = a2980 & ~a2020;
assign a2984 = a2982 & ~a2010;
assign a2986 = ~a2984 & ~a2008;
assign a2988 = ~a2986 & ~a2004;
assign a2990 = a2988 & ~a2000;
assign a2992 = a2990 & ~a1984;
assign a2994 = a2992 & ~a1980;
assign a2996 = a2994 & ~a1978;
assign a2998 = a2996 & ~a1976;
assign a3000 = a2998 & ~a1968;
assign a3002 = a3000 & ~a1966;
assign a3004 = a3002 & ~a1960;
assign a3006 = a3004 & ~a1950;
assign a3008 = a3006 & ~a1944;
assign a3010 = a3008 & ~a1938;
assign a3012 = a3010 & ~a1936;
assign a3014 = a3012 & ~a1934;
assign a3016 = a3014 & ~a1932;
assign a3018 = a3016 & ~a1930;
assign a3020 = ~a3018 & ~a1928;
assign a3022 = ~a3020 & ~a1916;
assign a3024 = a3022 & ~a1908;
assign a3026 = a3024 & ~a1892;
assign a3028 = a3026 & ~a1890;
assign a3030 = a3028 & ~a1884;
assign a3032 = a3030 & ~a1876;
assign a3034 = a3032 & ~a1866;
assign a3036 = a3034 & ~a1858;
assign a3038 = a3036 & ~a1850;
assign a3040 = a3038 & ~a1838;
assign a3042 = a3040 & ~a1834;
assign a3044 = a3042 & ~a1826;
assign a3046 = a3044 & ~a1824;
assign a3048 = a3046 & ~a1822;
assign a3050 = a3048 & ~a1820;
assign a3052 = a3050 & ~a1818;
assign a3054 = ~a3052 & ~a1810;
assign a3056 = ~a3054 & ~a1796;
assign a3058 = a3056 & ~a1786;
assign a3060 = a3058 & ~a1770;
assign a3062 = a3060 & ~a1768;
assign a3064 = a3062 & ~a1762;
assign a3066 = a3064 & ~a1754;
assign a3068 = a3066 & ~a1744;
assign a3070 = a3068 & ~a1736;
assign a3072 = a3070 & ~a1728;
assign a3074 = a3072 & ~a1716;
assign a3076 = a3074 & ~a1712;
assign a3078 = a3076 & ~a1704;
assign a3080 = a3078 & ~a1702;
assign a3082 = a3080 & ~a1700;
assign a3084 = a3082 & ~a1698;
assign a3086 = a3084 & ~a1696;
assign a3088 = ~a3086 & ~a1688;
assign a3090 = ~a3088 & ~a1674;
assign a3092 = a3090 & ~a1664;
assign a3094 = a3092 & ~a1648;
assign a3096 = a3094 & ~a1646;
assign a3098 = a3096 & ~a1640;
assign a3100 = a3098 & ~a1632;
assign a3102 = a3100 & ~a1624;
assign a3104 = a3102 & ~a1618;
assign a3106 = a3104 & ~a1606;
assign a3108 = a3106 & ~a1594;
assign a3110 = a3108 & ~a1590;
assign a3112 = a3110 & ~a1582;
assign a3114 = ~a3112 & ~a1574;
assign a3116 = a3114 & ~a1566;
assign a3118 = a3116 & ~a1558;
assign a3120 = ~a3118 & ~a1548;
assign a3122 = a3120 & ~a1538;
assign a3124 = a3122 & ~a1528;
assign a3126 = a3124 & ~a1522;
assign a3128 = a3126 & ~a1506;
assign a3130 = a3128 & ~a1502;
assign a3132 = a3130 & ~a1494;
assign a3134 = a3132 & ~a1486;
assign a3136 = a3134 & ~a1482;
assign a3138 = a3136 & ~a1478;
assign a3140 = a3138 & ~a1476;
assign a3142 = a3140 & ~a1472;
assign a3144 = a3142 & ~a1462;
assign a3146 = a3144 & ~a1448;
assign a3148 = a3146 & ~a1446;
assign a3150 = a3148 & ~a1442;
assign a3152 = a3150 & ~a1436;
assign a3154 = a3152 & ~a1428;
assign a3156 = a3154 & ~a1420;
assign a3158 = a3156 & ~a1418;
assign a3160 = a3158 & ~a1416;
assign a3162 = a3160 & ~a1414;
assign a3164 = ~a3162 & ~a1408;
assign a3166 = ~a3164 & ~a1404;
assign a3168 = a3166 & ~a1398;
assign a3170 = a3168 & ~a1392;
assign a3172 = a3170 & ~a1378;
assign a3174 = a3172 & ~a1376;
assign a3176 = a3174 & ~a1372;
assign a3178 = a3176 & ~a1364;
assign a3180 = a3178 & ~a1356;
assign a3182 = a3180 & ~a1352;
assign a3184 = a3182 & ~a1346;
assign a3186 = a3184 & ~a1338;
assign a3188 = a3186 & ~a1330;
assign a3190 = a3188 & ~a1320;
assign a3192 = a3190 & ~a1306;
assign a3194 = a3192 & ~a1290;
assign a3196 = a3194 & ~a1284;
assign a3198 = a3196 & ~a1278;
assign a3200 = a3198 & ~a1268;
assign a3202 = a3200 & ~a1254;
assign a3204 = a3202 & ~a1242;
assign a3206 = a3204 & ~a1230;
assign a3208 = a3206 & ~a1222;
assign a3210 = a3208 & ~a1214;
assign a3212 = a3210 & ~a1200;
assign a3214 = a3212 & ~a1198;
assign a3216 = a3214 & ~a1194;
assign a3218 = a3216 & ~a1186;
assign a3220 = a3218 & ~a1178;
assign a3222 = ~a3220 & ~a1176;
assign a3224 = ~a3222 & ~a1172;
assign a3226 = a3224 & ~a1162;
assign a3228 = a3226 & ~a1156;
assign a3230 = a3228 & ~a1152;
assign a3232 = a3230 & ~a1150;
assign a3234 = a3232 & ~a1140;
assign a3236 = a3234 & ~a1128;
assign a3238 = a3236 & ~a1116;
assign a3240 = a3238 & ~a1104;
assign a3242 = a3240 & ~a1100;
assign a3244 = a3242 & ~a1090;
assign a3246 = a3244 & ~a1080;
assign a3248 = a3246 & ~a1060;
assign a3250 = a3248 & ~a1056;
assign a3252 = a3250 & ~a1048;
assign a3254 = a3252 & ~a1040;
assign a3256 = a3254 & ~a1038;
assign a3258 = a3256 & ~a1032;
assign a3260 = a3258 & ~a1030;
assign a3262 = a3260 & ~a1024;
assign a3264 = a3262 & ~a1010;
assign a3266 = a3264 & ~a996;
assign a3268 = a3266 & ~a992;
assign a3270 = a3268 & ~a986;
assign a3272 = a3270 & ~a982;
assign a3274 = a3272 & ~a968;
assign a3276 = a3274 & ~a964;
assign a3278 = a3276 & ~a956;
assign a3280 = a3278 & ~a948;
assign a3282 = a3280 & ~a944;
assign a3284 = a3282 & ~a934;
assign a3286 = a3284 & ~a928;
assign a3288 = ~a3286 & ~a926;
assign a3290 = ~a3288 & ~a912;
assign a3292 = a3290 & ~a908;
assign a3294 = a3292 & ~a902;
assign a3296 = a3294 & ~a896;
assign a3298 = a3296 & ~a888;
assign a3300 = a3298 & ~a876;
assign a3302 = a3300 & ~a860;
assign a3304 = ~a3302 & i96;
assign a3306 = a3302 & ~i96;
assign a3308 = ~a3306 & ~a3304;
assign a3310 = a940 & l304;
assign a3312 = a3310 & l308;
assign a3314 = a3312 & ~l326;
assign a3316 = a920 & ~l304;
assign a3318 = a3316 & ~l326;
assign a3320 = a920 & ~l308;
assign a3322 = a3320 & ~l326;
assign a3324 = a972 & ~i106;
assign a3326 = a3324 & ~i110;
assign a3328 = a3326 & i108;
assign a3330 = a3328 & l304;
assign a3332 = a3330 & l326;
assign a3334 = a3328 & ~l304;
assign a3336 = a3334 & l326;
assign a3338 = a1694 & l302;
assign a3340 = a3338 & l304;
assign a3342 = a3340 & l308;
assign a3344 = a1682 & ~l302;
assign a3346 = a1682 & ~l304;
assign a3348 = a1682 & ~l308;
assign a3350 = a1730 & ~i106;
assign a3352 = a3350 & ~i110;
assign a3354 = a3352 & i108;
assign a3356 = a1816 & l302;
assign a3358 = a3356 & l304;
assign a3360 = a3358 & l308;
assign a3362 = a1804 & ~l302;
assign a3364 = a1804 & ~l304;
assign a3366 = a1804 & ~l308;
assign a3368 = a1852 & ~i106;
assign a3370 = a3368 & ~i110;
assign a3372 = a3370 & i108;
assign a3374 = a2044 & ~i106;
assign a3376 = a3374 & ~i110;
assign a3378 = a3376 & i108;
assign a3380 = a3378 & ~l304;
assign a3382 = a2266 & ~i106;
assign a3384 = a3382 & ~i110;
assign a3386 = a3384 & i108;
assign a3388 = a2334 & ~i106;
assign a3390 = a3388 & ~i110;
assign a3392 = a3390 & i108;
assign a3394 = a2440 & ~i106;
assign a3396 = a3394 & ~i110;
assign a3398 = a3396 & i108;
assign a3400 = a3398 & ~l326;
assign a3402 = a2496 & ~i106;
assign a3404 = a3402 & ~i110;
assign a3406 = a3404 & i108;
assign a3408 = a3406 & l326;
assign a3410 = a2588 & ~i106;
assign a3412 = a3410 & ~i110;
assign a3414 = a3412 & i108;
assign a3416 = a3414 & ~l326;
assign a3418 = a2660 & ~i106;
assign a3420 = a3418 & ~i110;
assign a3422 = a3420 & i108;
assign a3424 = a3422 & l326;
assign a3426 = a1066 & l268;
assign a3428 = a3426 & ~l236;
assign a3430 = a3428 & ~l294;
assign a3432 = a3430 & ~a1062;
assign a3434 = a3432 & i110;
assign a3436 = a3434 & ~i108;
assign a3438 = a3436 & i106;
assign a3440 = ~l274 & ~l270;
assign a3442 = a3440 & ~l236;
assign a3444 = l276 & ~l272;
assign a3446 = a3444 & l268;
assign a3448 = a3446 & ~a952;
assign a3450 = a3448 & i110;
assign a3452 = a3450 & i108;
assign a3454 = a3452 & ~i106;
assign a3456 = a3428 & ~a960;
assign a3458 = a3456 & i110;
assign a3460 = a3458 & ~i108;
assign a3462 = a3460 & ~i106;
assign a3464 = a3428 & ~l288;
assign a3466 = a3464 & l290;
assign a3468 = a3466 & ~i118;
assign a3470 = a3446 & l294;
assign a3472 = a3470 & ~a1062;
assign a3474 = a3472 & i110;
assign a3476 = a3474 & ~i108;
assign a3478 = a3476 & i106;
assign a3480 = a3464 & i116;
assign a3482 = ~l286 & l276;
assign a3484 = a3482 & i114;
assign a3486 = a3484 & l314;
assign a3488 = a2056 & ~l268;
assign a3490 = a3488 & ~l236;
assign a3492 = a3490 & i64;
assign a3494 = a3492 & ~l294;
assign a3496 = a3494 & l326;
assign a3498 = a3490 & ~l294;
assign a3500 = a3498 & ~a864;
assign a3502 = a3500 & ~i110;
assign a3504 = a3502 & i108;
assign a3506 = a3504 & ~i106;
assign a3508 = a3506 & l326;
assign a3510 = a3498 & ~a1062;
assign a3512 = a3510 & i110;
assign a3514 = a3512 & ~i108;
assign a3516 = a3514 & i106;
assign a3518 = a3516 & l326;
assign a3520 = ~a952 & l276;
assign a3522 = a3520 & i110;
assign a3524 = a3522 & i108;
assign a3526 = a3524 & ~i106;
assign a3528 = a3490 & ~a960;
assign a3530 = a3528 & i110;
assign a3532 = a3530 & ~i108;
assign a3534 = a3532 & ~i106;
assign a3536 = a3490 & ~l288;
assign a3538 = a3536 & l290;
assign a3540 = a3538 & ~i118;
assign a3542 = l294 & l276;
assign a3544 = a3542 & ~a864;
assign a3546 = a3544 & ~i106;
assign a3548 = a3546 & ~i110;
assign a3550 = a3548 & i108;
assign a3552 = a3550 & l326;
assign a3554 = a3536 & i116;
assign a3556 = a1062 & i64;
assign a3558 = a1082 & i64;
assign a3560 = ~l298 & i126;
assign a3562 = ~a3560 & ~i64;
assign a3564 = ~a3562 & a950;
assign a3566 = ~a3564 & ~a3558;
assign a3568 = ~a3566 & ~l278;
assign a3570 = a864 & i64;
assign a3572 = a1084 & l238;
assign a3574 = a3572 & ~l298;
assign a3576 = a3574 & i126;
assign a3578 = a864 & ~l298;
assign a3580 = a3578 & i126;
assign a3582 = a1062 & ~l298;
assign a3584 = a3582 & i126;
assign a3586 = a1084 & ~l238;
assign a3588 = a3586 & ~l298;
assign a3590 = a3588 & i126;
assign a3592 = ~a3590 & ~a3584;
assign a3594 = a3592 & ~a3580;
assign a3596 = a3594 & ~a3576;
assign a3598 = a3596 & ~a3570;
assign a3600 = a3598 & ~a3568;
assign a3602 = a3600 & ~a3556;
assign a3604 = l290 & ~l276;
assign a3606 = a3604 & ~a3602;
assign a3608 = a3606 & ~a3554;
assign a3610 = a3542 & ~a1062;
assign a3612 = a3610 & i110;
assign a3614 = a3612 & ~i108;
assign a3616 = a3614 & i106;
assign a3618 = a3616 & l326;
assign a3620 = l276 & i64;
assign a3622 = a3620 & l294;
assign a3624 = a3622 & l326;
assign a3626 = ~a3624 & ~a3618;
assign a3628 = a3626 & ~a3608;
assign a3630 = a3628 & ~a3552;
assign a3632 = ~a3630 & ~a3540;
assign a3634 = a3632 & ~a3534;
assign a3636 = l276 & l216;
assign a3638 = a3636 & ~i44;
assign a3640 = ~a864 & l276;
assign a3642 = a3640 & ~i106;
assign a3644 = a3642 & ~i110;
assign a3646 = a3644 & i108;
assign a3648 = a3646 & ~l326;
assign a3650 = a3648 & l330;
assign a3652 = ~a1062 & l276;
assign a3654 = a3652 & i110;
assign a3656 = a3654 & ~i108;
assign a3658 = a3656 & i106;
assign a3660 = a3658 & ~l326;
assign a3662 = a3660 & l330;
assign a3664 = a864 & l276;
assign a3666 = a3664 & ~l330;
assign a3668 = a3666 & i156;
assign a3670 = a1062 & l276;
assign a3672 = a3670 & ~l330;
assign a3674 = a3672 & i156;
assign a3676 = a3620 & a1084;
assign a3678 = a3676 & ~l326;
assign a3680 = a3620 & a1062;
assign a3682 = a3620 & a864;
assign a3684 = ~a3682 & ~a3680;
assign a3686 = a3684 & ~a3678;
assign a3688 = a3686 & ~a3674;
assign a3690 = a3688 & ~a3668;
assign a3692 = a3690 & ~a3662;
assign a3694 = a3692 & ~a3650;
assign a3696 = a3694 & ~a3638;
assign a3698 = a3696 & ~a3634;
assign a3700 = a3698 & ~a3526;
assign a3702 = ~a3700 & ~a3518;
assign a3704 = a3702 & ~a3508;
assign a3706 = a3704 & ~a3496;
assign a3708 = ~a3706 & ~a3486;
assign a3710 = l272 & ~l268;
assign a3712 = a3710 & ~a3708;
assign a3714 = a3712 & ~a3480;
assign a3716 = a3470 & ~a864;
assign a3718 = a3716 & ~i106;
assign a3720 = a3718 & ~i110;
assign a3722 = a3720 & i108;
assign a3724 = a3446 & i64;
assign a3726 = a3724 & l294;
assign a3728 = ~a3726 & ~a3722;
assign a3730 = a3728 & ~a3714;
assign a3732 = a3730 & ~a3478;
assign a3734 = ~a3732 & ~a3468;
assign a3736 = a3734 & ~a3462;
assign a3738 = ~a3736 & ~a3454;
assign a3740 = a3430 & ~a864;
assign a3742 = a3740 & ~i110;
assign a3744 = a3742 & i108;
assign a3746 = a3744 & ~i106;
assign a3748 = a3428 & i64;
assign a3750 = a3748 & ~l294;
assign a3752 = a3428 & ~l216;
assign a3754 = a3752 & i44;
assign a3756 = ~a3754 & ~a3750;
assign a3758 = a3756 & ~a3746;
assign a3760 = a3758 & ~a3738;
assign a3762 = a3760 & a3442;
assign a3764 = a3762 & ~a3438;
assign a3766 = ~a3764 & ~l270;
assign a3768 = a3766 & ~a2694;
assign a3770 = a3768 & ~a2688;
assign a3772 = ~a3770 & ~a2680;
assign a3774 = ~a3772 & ~a2678;
assign a3776 = a3774 & ~a3424;
assign a3778 = a3776 & ~a2656;
assign a3780 = a3778 & ~a2644;
assign a3782 = ~a3780 & ~a2640;
assign a3784 = a3782 & ~a2634;
assign a3786 = ~a3784 & ~a2626;
assign a3788 = a3786 & ~a2618;
assign a3790 = a3788 & ~a2616;
assign a3792 = a3790 & ~a2606;
assign a3794 = a3792 & ~a3416;
assign a3796 = ~a3794 & ~a2586;
assign a3798 = a3796 & ~a2576;
assign a3800 = a3798 & ~a2564;
assign a3802 = a3800 & ~a2550;
assign a3804 = ~a3802 & ~a2544;
assign a3806 = a3804 & ~a2538;
assign a3808 = a3806 & ~a2532;
assign a3810 = ~a3808 & ~a2516;
assign a3812 = ~a3810 & ~a2514;
assign a3814 = a3812 & ~a3408;
assign a3816 = a3814 & ~a2492;
assign a3818 = a3816 & ~a2488;
assign a3820 = ~a3818 & ~a2484;
assign a3822 = a3820 & ~a2478;
assign a3824 = ~a3822 & ~a2470;
assign a3826 = a3824 & ~a2462;
assign a3828 = a3826 & ~a2460;
assign a3830 = a3828 & ~a2458;
assign a3832 = a3830 & ~a3400;
assign a3834 = ~a3832 & ~a2438;
assign a3836 = a3834 & ~a2428;
assign a3838 = a3836 & ~a2416;
assign a3840 = a3838 & ~a2408;
assign a3842 = a3840 & ~a2402;
assign a3844 = ~a3842 & ~a2398;
assign a3846 = a3844 & ~a2392;
assign a3848 = ~a3846 & ~a2380;
assign a3850 = ~a3848 & ~a2378;
assign a3852 = ~a3850 & ~a2372;
assign a3854 = a3852 & ~a2368;
assign a3856 = ~a3854 & ~a2360;
assign a3858 = a3856 & ~a2352;
assign a3860 = a3858 & ~a2342;
assign a3862 = a3860 & ~a3392;
assign a3864 = a3862 & ~a2332;
assign a3866 = ~a3864 & ~a2324;
assign a3868 = ~a3866 & ~a2314;
assign a3870 = ~a3868 & ~a2302;
assign a3872 = ~a3870 & ~a2300;
assign a3874 = ~a3872 & ~a2294;
assign a3876 = a3874 & ~a2290;
assign a3878 = ~a3876 & ~a2282;
assign a3880 = a3878 & ~a2274;
assign a3882 = a3880 & ~a3386;
assign a3884 = a3882 & ~a2264;
assign a3886 = ~a3884 & ~a2256;
assign a3888 = ~a3886 & ~a2246;
assign a3890 = ~a3888 & ~a2234;
assign a3892 = a3890 & ~a2232;
assign a3894 = a3892 & ~a2226;
assign a3896 = ~a3894 & ~a2218;
assign a3898 = a3896 & ~a2210;
assign a3900 = a3898 & ~a2208;
assign a3902 = a3900 & ~a2206;
assign a3904 = ~a3902 & ~a2204;
assign a3906 = a3904 & ~a2198;
assign a3908 = ~a3906 & ~a2194;
assign a3910 = a3908 & ~a2188;
assign a3912 = a3910 & ~a2182;
assign a3914 = a3912 & ~a2168;
assign a3916 = a3914 & ~a2166;
assign a3918 = a3916 & ~a2164;
assign a3920 = a3918 & ~a2158;
assign a3922 = a3920 & ~a2156;
assign a3924 = a3922 & ~a2154;
assign a3926 = ~a3924 & ~a2146;
assign a3928 = a3926 & ~a2142;
assign a3930 = ~a3928 & ~a2134;
assign a3932 = a3930 & ~a2126;
assign a3934 = a3932 & ~a2124;
assign a3936 = ~a3934 & ~a2122;
assign a3938 = a3936 & ~a2118;
assign a3940 = a3938 & ~a2108;
assign a3942 = a3940 & ~a2096;
assign a3944 = a3942 & ~a2084;
assign a3946 = a3944 & ~a2076;
assign a3948 = ~a3946 & ~a2068;
assign a3950 = a3948 & ~a2054;
assign a3952 = a3950 & ~a3380;
assign a3954 = a3952 & ~a2042;
assign a3956 = a3954 & ~a2036;
assign a3958 = ~a3956 & ~a2032;
assign a3960 = a3958 & ~a2028;
assign a3962 = ~a3960 & ~a2020;
assign a3964 = a3962 & ~a2010;
assign a3966 = ~a3964 & ~a2008;
assign a3968 = a3966 & ~a2004;
assign a3970 = a3968 & ~a2000;
assign a3972 = a3970 & ~a1984;
assign a3974 = a3972 & ~a1980;
assign a3976 = ~a3974 & ~a1978;
assign a3978 = a3976 & ~a1976;
assign a3980 = a3978 & ~a1968;
assign a3982 = a3980 & ~a1966;
assign a3984 = a3982 & ~a1960;
assign a3986 = ~a3984 & ~a1950;
assign a3988 = ~a3986 & ~a1944;
assign a3990 = a3988 & ~a1938;
assign a3992 = a3990 & ~a1936;
assign a3994 = a3992 & ~a1934;
assign a3996 = a3994 & ~a1932;
assign a3998 = a3996 & ~a1930;
assign a4000 = ~a3998 & ~a1928;
assign a4002 = a4000 & ~a1916;
assign a4004 = a4002 & ~a1908;
assign a4006 = a4004 & ~a1892;
assign a4008 = a4006 & ~a1890;
assign a4010 = ~a4008 & ~a1884;
assign a4012 = a4010 & ~a1876;
assign a4014 = a4012 & ~a1866;
assign a4016 = a4014 & ~a3372;
assign a4018 = a4016 & ~a1850;
assign a4020 = ~a4018 & ~a1838;
assign a4022 = ~a4020 & ~a1834;
assign a4024 = a4022 & ~a1826;
assign a4026 = a4024 & ~a1824;
assign a4028 = a4026 & ~a3366;
assign a4030 = a4028 & ~a3364;
assign a4032 = a4030 & ~a3362;
assign a4034 = ~a4032 & ~a3360;
assign a4036 = a4034 & ~a1796;
assign a4038 = a4036 & ~a1786;
assign a4040 = a4038 & ~a1770;
assign a4042 = a4040 & ~a1768;
assign a4044 = a4042 & ~a1762;
assign a4046 = ~a4044 & ~a1754;
assign a4048 = a4046 & ~a1744;
assign a4050 = a4048 & ~a3354;
assign a4052 = a4050 & ~a1728;
assign a4054 = ~a4052 & ~a1716;
assign a4056 = a4054 & ~a1712;
assign a4058 = ~a4056 & ~a1704;
assign a4060 = a4058 & ~a1702;
assign a4062 = a4060 & ~a3348;
assign a4064 = a4062 & ~a3346;
assign a4066 = a4064 & ~a3344;
assign a4068 = ~a4066 & ~a3342;
assign a4070 = a4068 & ~a1674;
assign a4072 = a4070 & ~a1664;
assign a4074 = a4072 & ~a1648;
assign a4076 = a4074 & ~a1646;
assign a4078 = a4076 & ~a1640;
assign a4080 = ~a4078 & ~a1632;
assign a4082 = ~a4080 & ~a1624;
assign a4084 = ~a4082 & ~a1618;
assign a4086 = a4084 & ~a1606;
assign a4088 = ~a4086 & ~a1594;
assign a4090 = a4088 & ~a1590;
assign a4092 = ~a4090 & ~a1582;
assign a4094 = ~a4092 & ~a1574;
assign a4096 = a4094 & ~a1566;
assign a4098 = a4096 & ~a1558;
assign a4100 = a4098 & ~a1548;
assign a4102 = a4100 & ~a1538;
assign a4104 = a4102 & ~a1528;
assign a4106 = a4104 & ~a1522;
assign a4108 = a4106 & ~a1506;
assign a4110 = a4108 & ~a1502;
assign a4112 = ~a4110 & ~a1494;
assign a4114 = a4112 & ~a1486;
assign a4116 = a4114 & ~a1482;
assign a4118 = a4116 & ~a1478;
assign a4120 = a4118 & ~a1476;
assign a4122 = ~a4120 & ~a1472;
assign a4124 = a4122 & ~a1462;
assign a4126 = a4124 & ~a1448;
assign a4128 = ~a4126 & ~a1446;
assign a4130 = ~a4128 & ~a1442;
assign a4132 = a4130 & ~a1436;
assign a4134 = ~a4132 & ~a1428;
assign a4136 = a4134 & ~a1420;
assign a4138 = a4136 & ~a1418;
assign a4140 = a4138 & ~a1416;
assign a4142 = ~a4140 & ~a1414;
assign a4144 = a4142 & ~a1408;
assign a4146 = ~a4144 & ~a1404;
assign a4148 = a4146 & ~a1398;
assign a4150 = a4148 & ~a1392;
assign a4152 = a4150 & ~a1378;
assign a4154 = ~a4152 & ~a1376;
assign a4156 = a4154 & ~a1372;
assign a4158 = ~a4156 & ~a1364;
assign a4160 = a4158 & ~a1356;
assign a4162 = ~a4160 & ~a1352;
assign a4164 = a4162 & ~a1346;
assign a4166 = a4164 & ~a1338;
assign a4168 = a4166 & ~a1330;
assign a4170 = a4168 & ~a1320;
assign a4172 = a4170 & ~a1306;
assign a4174 = a4172 & ~a1290;
assign a4176 = a4174 & ~a1284;
assign a4178 = a4176 & ~a1278;
assign a4180 = a4178 & ~a1268;
assign a4182 = a4180 & ~a1254;
assign a4184 = a4182 & ~a1242;
assign a4186 = a4184 & ~a1230;
assign a4188 = a4186 & ~a1222;
assign a4190 = ~a4188 & ~a1214;
assign a4192 = a4190 & ~a1200;
assign a4194 = ~a4192 & ~a1198;
assign a4196 = a4194 & ~a1194;
assign a4198 = ~a4196 & ~a1186;
assign a4200 = a4198 & ~a1178;
assign a4202 = ~a4200 & ~a1176;
assign a4204 = a4202 & ~a1172;
assign a4206 = a4204 & ~a1162;
assign a4208 = a4206 & ~a1156;
assign a4210 = a4208 & ~a1152;
assign a4212 = a4210 & ~a1150;
assign a4214 = a4212 & ~a1140;
assign a4216 = a4214 & ~a1128;
assign a4218 = a4216 & ~a1116;
assign a4220 = a4218 & ~a1104;
assign a4222 = a4220 & ~a1100;
assign a4224 = a4222 & ~a1090;
assign a4226 = a4224 & ~a1080;
assign a4228 = a4226 & ~a1060;
assign a4230 = a4228 & ~a1056;
assign a4232 = ~a4230 & ~a1048;
assign a4234 = ~a4232 & ~a1040;
assign a4236 = a4234 & ~a1038;
assign a4238 = a4236 & ~a1032;
assign a4240 = a4238 & ~a1030;
assign a4242 = a4240 & ~a1024;
assign a4244 = a4242 & ~a1010;
assign a4246 = ~a4244 & ~a3336;
assign a4248 = a4246 & ~a992;
assign a4250 = a4248 & ~a986;
assign a4252 = a4250 & ~a3332;
assign a4254 = ~a4252 & ~a968;
assign a4256 = a4254 & ~a964;
assign a4258 = ~a4256 & ~a956;
assign a4260 = a4258 & ~a3322;
assign a4262 = a4260 & ~a3318;
assign a4264 = a4262 & ~a934;
assign a4266 = a4264 & ~a928;
assign a4268 = ~a4266 & ~a3314;
assign a4270 = a4268 & ~a912;
assign a4272 = a4270 & ~a908;
assign a4274 = a4272 & ~a902;
assign a4276 = a4274 & ~a896;
assign a4278 = a4276 & ~a888;
assign a4280 = a4278 & ~a876;
assign a4282 = a4280 & ~a860;
assign a4284 = ~a4282 & i98;
assign a4286 = a4282 & ~i98;
assign a4288 = ~a4286 & ~a4284;
assign a4290 = ~i110 & ~i106;
assign a4292 = a4290 & i108;
assign a4294 = a4292 & a890;
assign a4296 = a4294 & ~l304;
assign a4298 = a4296 & l326;
assign a4300 = a1014 & ~i106;
assign a4302 = a4300 & ~i110;
assign a4304 = a4302 & i108;
assign a4306 = a4304 & ~l304;
assign a4308 = a1164 & ~i106;
assign a4310 = a4308 & ~i110;
assign a4312 = a4310 & i108;
assign a4314 = a4312 & ~l304;
assign a4316 = a2420 & ~i106;
assign a4318 = a4316 & ~i110;
assign a4320 = a4318 & i108;
assign a4322 = a4320 & l326;
assign a4324 = a2568 & ~i106;
assign a4326 = a4324 & ~i110;
assign a4328 = a4326 & i108;
assign a4330 = a4328 & l326;
assign a4332 = a2706 & ~i106;
assign a4334 = a4332 & ~i110;
assign a4336 = a4334 & i108;
assign a4338 = a2748 & ~i106;
assign a4340 = a4338 & ~i110;
assign a4342 = a4340 & i108;
assign a4344 = a2056 & ~l270;
assign a4346 = a4344 & ~l268;
assign a4348 = a4346 & ~l236;
assign a4350 = a4348 & ~l286;
assign a4352 = a4350 & i114;
assign a4354 = a4352 & l314;
assign a4356 = a1064 & ~l270;
assign a4358 = a4356 & ~l268;
assign a4360 = a4358 & ~l236;
assign a4362 = a4360 & ~l294;
assign a4364 = a4362 & ~a1062;
assign a4366 = a4364 & i110;
assign a4368 = a4366 & ~i108;
assign a4370 = a4368 & i106;
assign a4372 = a4370 & l326;
assign a4374 = ~l274 & l272;
assign a4376 = a4374 & ~l270;
assign a4378 = a4376 & ~l268;
assign a4380 = a4378 & ~l236;
assign a4382 = ~a960 & l276;
assign a4384 = a4382 & i110;
assign a4386 = a4384 & ~i108;
assign a4388 = a4386 & ~i106;
assign a4390 = a4360 & ~l288;
assign a4392 = a4390 & l290;
assign a4394 = a4392 & ~i118;
assign a4396 = a4360 & i64;
assign a4398 = a4396 & l294;
assign a4400 = a4398 & l326;
assign a4402 = a4360 & l294;
assign a4404 = a4402 & ~a1062;
assign a4406 = a4404 & i110;
assign a4408 = a4406 & ~i108;
assign a4410 = a4408 & i106;
assign a4412 = a4410 & l326;
assign a4414 = a4402 & ~a864;
assign a4416 = a4414 & ~i106;
assign a4418 = a4416 & ~i110;
assign a4420 = a4418 & i108;
assign a4422 = a4420 & l326;
assign a4424 = a4390 & i116;
assign a4426 = l280 & i64;
assign a4428 = ~a3562 & ~l280;
assign a4430 = ~l298 & l280;
assign a4432 = a4430 & i126;
assign a4434 = ~a4432 & ~a4428;
assign a4436 = a4434 & ~a4426;
assign a4438 = ~a4436 & l282;
assign a4440 = ~a4438 & ~a3558;
assign a4442 = ~a4440 & ~l278;
assign a4444 = ~a4442 & a3598;
assign a4446 = a4444 & ~a3556;
assign a4448 = ~a4446 & a3604;
assign a4450 = a4448 & ~a4424;
assign a4452 = a4450 & ~a4422;
assign a4454 = a4452 & ~a4412;
assign a4456 = a4454 & ~a4400;
assign a4458 = a4456 & ~a4394;
assign a4460 = a3640 & ~i110;
assign a4462 = a4460 & i108;
assign a4464 = a4462 & ~i106;
assign a4466 = a4464 & ~l326;
assign a4468 = a4466 & l330;
assign a4470 = ~a4468 & a3692;
assign a4472 = a4470 & ~a3638;
assign a4474 = a4472 & ~a3526;
assign a4476 = a4474 & ~a4458;
assign a4478 = a4476 & ~a4388;
assign a4480 = a4362 & ~a864;
assign a4482 = a4480 & ~i106;
assign a4484 = a4482 & ~i110;
assign a4486 = a4484 & i108;
assign a4488 = a4486 & l326;
assign a4490 = a4396 & ~l294;
assign a4492 = a4490 & l326;
assign a4494 = ~a4492 & ~a4488;
assign a4496 = a4494 & ~a4478;
assign a4498 = a4496 & a4380;
assign a4500 = a4498 & ~a4372;
assign a4502 = ~a4500 & l272;
assign a4504 = a4502 & ~a4354;
assign a4506 = ~a4504 & ~a2764;
assign a4508 = a4506 & ~a2762;
assign a4510 = a4508 & ~a4342;
assign a4512 = a4510 & ~a2744;
assign a4514 = a4512 & ~a2742;
assign a4516 = ~a4514 & ~a2736;
assign a4518 = a4516 & ~a2728;
assign a4520 = ~a4518 & ~a2720;
assign a4522 = a4520 & ~a4336;
assign a4524 = a4522 & ~a2702;
assign a4526 = a4524 & ~a2698;
assign a4528 = ~a4526 & ~a2694;
assign a4530 = a4528 & ~a2688;
assign a4532 = ~a4530 & ~a2680;
assign a4534 = a4532 & ~a2678;
assign a4536 = a4534 & ~a3424;
assign a4538 = a4536 & ~a2656;
assign a4540 = a4538 & ~a2644;
assign a4542 = a4540 & ~a2640;
assign a4544 = ~a4542 & ~a2634;
assign a4546 = a4544 & ~a2626;
assign a4548 = a4546 & ~a2618;
assign a4550 = a4548 & ~a2616;
assign a4552 = a4550 & ~a2606;
assign a4554 = a4552 & ~a2596;
assign a4556 = ~a4554 & ~a2586;
assign a4558 = a4556 & ~a4330;
assign a4560 = a4558 & ~a2564;
assign a4562 = a4560 & ~a2550;
assign a4564 = a4562 & ~a2544;
assign a4566 = ~a4564 & ~a2538;
assign a4568 = ~a4566 & ~a2532;
assign a4570 = a4568 & ~a2516;
assign a4572 = a4570 & ~a2514;
assign a4574 = a4572 & ~a3408;
assign a4576 = a4574 & ~a2492;
assign a4578 = a4576 & ~a2488;
assign a4580 = a4578 & ~a2484;
assign a4582 = ~a4580 & ~a2478;
assign a4584 = a4582 & ~a2470;
assign a4586 = a4584 & ~a2462;
assign a4588 = a4586 & ~a2460;
assign a4590 = a4588 & ~a2458;
assign a4592 = a4590 & ~a2448;
assign a4594 = ~a4592 & ~a2438;
assign a4596 = a4594 & ~a4322;
assign a4598 = a4596 & ~a2416;
assign a4600 = a4598 & ~a2408;
assign a4602 = a4600 & ~a2402;
assign a4604 = ~a4602 & ~a2398;
assign a4606 = a4604 & ~a2392;
assign a4608 = ~a4606 & ~a2380;
assign a4610 = a4608 & ~a2378;
assign a4612 = a4610 & ~a2372;
assign a4614 = ~a4612 & ~a2368;
assign a4616 = a4614 & ~a2360;
assign a4618 = a4616 & ~a2352;
assign a4620 = a4618 & ~a2342;
assign a4622 = a4620 & ~a2340;
assign a4624 = a4622 & ~a2332;
assign a4626 = ~a4624 & ~a2324;
assign a4628 = a4626 & ~a2314;
assign a4630 = a4628 & ~a2302;
assign a4632 = a4630 & ~a2300;
assign a4634 = a4632 & ~a2294;
assign a4636 = ~a4634 & ~a2290;
assign a4638 = a4636 & ~a2282;
assign a4640 = a4638 & ~a2274;
assign a4642 = a4640 & ~a2272;
assign a4644 = a4642 & ~a2264;
assign a4646 = ~a4644 & ~a2256;
assign a4648 = ~a4646 & ~a2246;
assign a4650 = ~a4648 & ~a2234;
assign a4652 = a4650 & ~a2232;
assign a4654 = ~a4652 & ~a2226;
assign a4656 = a4654 & ~a2218;
assign a4658 = a4656 & ~a2210;
assign a4660 = a4658 & ~a2208;
assign a4662 = a4660 & ~a2206;
assign a4664 = ~a4662 & ~a2204;
assign a4666 = ~a4664 & ~a2198;
assign a4668 = ~a4666 & ~a2194;
assign a4670 = ~a4668 & ~a2188;
assign a4672 = a4670 & ~a2182;
assign a4674 = ~a4672 & ~a2168;
assign a4676 = a4674 & ~a2166;
assign a4678 = a4676 & ~a2164;
assign a4680 = a4678 & ~a2158;
assign a4682 = a4680 & ~a2156;
assign a4684 = a4682 & ~a2154;
assign a4686 = a4684 & ~a2146;
assign a4688 = ~a4686 & ~a2142;
assign a4690 = a4688 & ~a2134;
assign a4692 = a4690 & ~a2126;
assign a4694 = a4692 & ~a2124;
assign a4696 = a4694 & ~a2122;
assign a4698 = a4696 & ~a2118;
assign a4700 = a4698 & ~a2108;
assign a4702 = a4700 & ~a2096;
assign a4704 = a4702 & ~a2084;
assign a4706 = a4704 & ~a2076;
assign a4708 = a4706 & ~a2068;
assign a4710 = ~a4708 & ~a2054;
assign a4712 = a4710 & ~a3380;
assign a4714 = a4712 & ~a2042;
assign a4716 = a4714 & ~a2036;
assign a4718 = a4716 & ~a2032;
assign a4720 = ~a4718 & ~a2028;
assign a4722 = a4720 & ~a2020;
assign a4724 = a4722 & ~a2010;
assign a4726 = a4724 & ~a2008;
assign a4728 = a4726 & ~a2004;
assign a4730 = a4728 & ~a2000;
assign a4732 = ~a4730 & ~a1984;
assign a4734 = ~a4732 & ~a1980;
assign a4736 = a4734 & ~a1978;
assign a4738 = a4736 & ~a1976;
assign a4740 = a4738 & ~a1968;
assign a4742 = a4740 & ~a1966;
assign a4744 = a4742 & ~a1960;
assign a4746 = a4744 & ~a1950;
assign a4748 = a4746 & ~a1944;
assign a4750 = a4748 & ~a1938;
assign a4752 = a4750 & ~a1936;
assign a4754 = a4752 & ~a1934;
assign a4756 = a4754 & ~a1932;
assign a4758 = a4756 & ~a1930;
assign a4760 = a4758 & ~a1928;
assign a4762 = a4760 & ~a1916;
assign a4764 = a4762 & ~a1908;
assign a4766 = ~a4764 & ~a1892;
assign a4768 = a4766 & ~a1890;
assign a4770 = ~a4768 & ~a1884;
assign a4772 = a4770 & ~a1876;
assign a4774 = a4772 & ~a1866;
assign a4776 = a4774 & ~a1858;
assign a4778 = a4776 & ~a1850;
assign a4780 = ~a4778 & ~a1838;
assign a4782 = ~a4780 & ~a1834;
assign a4784 = a4782 & ~a1826;
assign a4786 = a4784 & ~a1824;
assign a4788 = a4786 & ~a1822;
assign a4790 = a4788 & ~a1820;
assign a4792 = a4790 & ~a1818;
assign a4794 = a4792 & ~a3360;
assign a4796 = a4794 & ~a1796;
assign a4798 = a4796 & ~a1786;
assign a4800 = ~a4798 & ~a1770;
assign a4802 = a4800 & ~a1768;
assign a4804 = ~a4802 & ~a1762;
assign a4806 = a4804 & ~a1754;
assign a4808 = a4806 & ~a1744;
assign a4810 = a4808 & ~a1736;
assign a4812 = a4810 & ~a1728;
assign a4814 = ~a4812 & ~a1716;
assign a4816 = ~a4814 & ~a1712;
assign a4818 = a4816 & ~a1704;
assign a4820 = a4818 & ~a1702;
assign a4822 = a4820 & ~a1700;
assign a4824 = a4822 & ~a1698;
assign a4826 = a4824 & ~a1696;
assign a4828 = a4826 & ~a3342;
assign a4830 = a4828 & ~a1674;
assign a4832 = a4830 & ~a1664;
assign a4834 = ~a4832 & ~a1648;
assign a4836 = a4834 & ~a1646;
assign a4838 = ~a4836 & ~a1640;
assign a4840 = a4838 & ~a1632;
assign a4842 = ~a4840 & ~a1624;
assign a4844 = a4842 & ~a1618;
assign a4846 = ~a4844 & ~a1606;
assign a4848 = ~a4846 & ~a1594;
assign a4850 = ~a4848 & ~a1590;
assign a4852 = a4850 & ~a1582;
assign a4854 = a4852 & ~a1574;
assign a4856 = a4854 & ~a1566;
assign a4858 = a4856 & ~a1558;
assign a4860 = a4858 & ~a1548;
assign a4862 = a4860 & ~a1538;
assign a4864 = a4862 & ~a1528;
assign a4866 = a4864 & ~a1522;
assign a4868 = ~a4866 & ~a1506;
assign a4870 = ~a4868 & ~a1502;
assign a4872 = a4870 & ~a1494;
assign a4874 = a4872 & ~a1486;
assign a4876 = a4874 & ~a1482;
assign a4878 = a4876 & ~a1478;
assign a4880 = a4878 & ~a1476;
assign a4882 = a4880 & ~a1472;
assign a4884 = a4882 & ~a1462;
assign a4886 = ~a4884 & ~a1448;
assign a4888 = a4886 & ~a1446;
assign a4890 = a4888 & ~a1442;
assign a4892 = ~a4890 & ~a1436;
assign a4894 = a4892 & ~a1428;
assign a4896 = a4894 & ~a1420;
assign a4898 = a4896 & ~a1418;
assign a4900 = a4898 & ~a1416;
assign a4902 = ~a4900 & ~a1414;
assign a4904 = ~a4902 & ~a1408;
assign a4906 = ~a4904 & ~a1404;
assign a4908 = ~a4906 & ~a1398;
assign a4910 = a4908 & ~a1392;
assign a4912 = ~a4910 & ~a1378;
assign a4914 = a4912 & ~a1376;
assign a4916 = ~a4914 & ~a1372;
assign a4918 = a4916 & ~a1364;
assign a4920 = a4918 & ~a1356;
assign a4922 = a4920 & ~a1352;
assign a4924 = a4922 & ~a1346;
assign a4926 = a4924 & ~a1338;
assign a4928 = a4926 & ~a1330;
assign a4930 = a4928 & ~a1320;
assign a4932 = a4930 & ~a1306;
assign a4934 = a4932 & ~a1290;
assign a4936 = a4934 & ~a1284;
assign a4938 = a4936 & ~a1278;
assign a4940 = a4938 & ~a1268;
assign a4942 = a4940 & ~a1254;
assign a4944 = a4942 & ~a1242;
assign a4946 = a4944 & ~a1230;
assign a4948 = a4946 & ~a1222;
assign a4950 = a4948 & ~a1214;
assign a4952 = ~a4950 & ~a1200;
assign a4954 = a4952 & ~a1198;
assign a4956 = ~a4954 & ~a1194;
assign a4958 = a4956 & ~a1186;
assign a4960 = a4958 & ~a1178;
assign a4962 = a4960 & ~a1176;
assign a4964 = ~a4962 & ~a4314;
assign a4966 = a4964 & ~a1162;
assign a4968 = a4966 & ~a1156;
assign a4970 = a4968 & ~a1152;
assign a4972 = ~a4970 & ~a1150;
assign a4974 = a4972 & ~a1140;
assign a4976 = a4974 & ~a1128;
assign a4978 = a4976 & ~a1116;
assign a4980 = a4978 & ~a1104;
assign a4982 = a4980 & ~a1100;
assign a4984 = a4982 & ~a1090;
assign a4986 = a4984 & ~a1080;
assign a4988 = ~a4986 & ~a1060;
assign a4990 = ~a4988 & ~a1056;
assign a4992 = a4990 & ~a1048;
assign a4994 = ~a4992 & ~a4306;
assign a4996 = a4994 & ~a1038;
assign a4998 = a4996 & ~a1032;
assign a5000 = ~a4998 & ~a1030;
assign a5002 = a5000 & ~a1024;
assign a5004 = a5002 & ~a1010;
assign a5006 = ~a5004 & ~a3336;
assign a5008 = a5006 & ~a992;
assign a5010 = a5008 & ~a986;
assign a5012 = a5010 & ~a3332;
assign a5014 = a5012 & ~a968;
assign a5016 = ~a5014 & ~a964;
assign a5018 = a5016 & ~a956;
assign a5020 = a5018 & ~a948;
assign a5022 = a5020 & ~a944;
assign a5024 = a5022 & ~a934;
assign a5026 = a5024 & ~a928;
assign a5028 = a5026 & ~a3314;
assign a5030 = ~a5028 & ~a4298;
assign a5032 = a5030 & ~a908;
assign a5034 = a5032 & ~a902;
assign a5036 = ~a5034 & ~a896;
assign a5038 = a5036 & ~a888;
assign a5040 = a5038 & ~a876;
assign a5042 = a5040 & ~a860;
assign a5044 = ~a5042 & i100;
assign a5046 = a5042 & ~i100;
assign a5048 = ~a5046 & ~a5044;
assign a5050 = a3444 & ~l270;
assign a5052 = a5050 & l268;
assign a5054 = a5052 & ~l236;
assign a5056 = a5054 & ~l216;
assign a5058 = a5056 & i44;
assign a5060 = a3446 & ~l288;
assign a5062 = a5060 & l290;
assign a5064 = a5062 & ~i118;
assign a5066 = a5054 & i64;
assign a5068 = a5066 & l294;
assign a5070 = a5054 & l294;
assign a5072 = a5070 & ~a864;
assign a5074 = a5072 & ~i110;
assign a5076 = a5074 & i108;
assign a5078 = a5076 & ~i106;
assign a5080 = a5070 & ~a1062;
assign a5082 = a5080 & i110;
assign a5084 = a5082 & ~i108;
assign a5086 = a5084 & i106;
assign a5088 = a5054 & ~l288;
assign a5090 = a5088 & i116;
assign a5092 = l276 & l272;
assign a5094 = a5092 & ~l270;
assign a5096 = a5094 & ~l268;
assign a5098 = a5096 & ~l236;
assign a5100 = a5098 & ~l286;
assign a5102 = a5100 & i114;
assign a5104 = a5102 & l314;
assign a5106 = ~l288 & l276;
assign a5108 = a5106 & l290;
assign a5110 = a5108 & ~i118;
assign a5112 = a5098 & i64;
assign a5114 = a5112 & l294;
assign a5116 = a5114 & l326;
assign a5118 = a5098 & l294;
assign a5120 = a5118 & ~a1062;
assign a5122 = a5120 & i110;
assign a5124 = a5122 & ~i108;
assign a5126 = a5124 & i106;
assign a5128 = a5126 & l326;
assign a5130 = a5118 & ~a864;
assign a5132 = a5130 & ~i110;
assign a5134 = a5132 & i108;
assign a5136 = a5134 & ~i106;
assign a5138 = a5136 & l326;
assign a5140 = a5098 & ~l288;
assign a5142 = a5140 & i116;
assign a5144 = ~l276 & l272;
assign a5146 = a5144 & ~l270;
assign a5148 = a5146 & ~l268;
assign a5150 = a5148 & ~l236;
assign a5152 = a5150 & ~l238;
assign a5154 = a5152 & l290;
assign a5156 = a5154 & a1084;
assign a5158 = a5156 & ~l298;
assign a5160 = a5158 & i126;
assign a5162 = l290 & i64;
assign a5164 = a5162 & a960;
assign a5166 = ~a3562 & ~l290;
assign a5168 = a960 & l290;
assign a5170 = a5168 & ~l298;
assign a5172 = a5170 & i126;
assign a5174 = a5162 & a952;
assign a5176 = a952 & l290;
assign a5178 = a5176 & ~l298;
assign a5180 = a5178 & i126;
assign a5182 = a5162 & a1084;
assign a5184 = a5162 & a1062;
assign a5186 = a5162 & a864;
assign a5188 = l290 & l238;
assign a5190 = a5188 & a1084;
assign a5192 = a5190 & ~l298;
assign a5194 = a5192 & i126;
assign a5196 = a864 & l290;
assign a5198 = a5196 & ~l298;
assign a5200 = a5198 & i126;
assign a5202 = a1062 & l290;
assign a5204 = a5202 & ~l298;
assign a5206 = a5204 & i126;
assign a5208 = ~a5206 & ~a5200;
assign a5210 = a5208 & ~a5194;
assign a5212 = a5210 & ~a5186;
assign a5214 = a5212 & ~a5184;
assign a5216 = a5214 & ~a5182;
assign a5218 = a5216 & ~a5180;
assign a5220 = a5218 & ~a5174;
assign a5222 = a5220 & ~a5172;
assign a5224 = a5222 & ~a5166;
assign a5226 = a5224 & ~a5164;
assign a5228 = ~a5226 & ~l276;
assign a5230 = a5228 & ~a5160;
assign a5232 = a5230 & ~a5142;
assign a5234 = a5232 & ~a5138;
assign a5236 = a5234 & ~a5128;
assign a5238 = a5236 & ~a5116;
assign a5240 = ~l294 & l276;
assign a5242 = a5240 & ~a1062;
assign a5244 = a5242 & i110;
assign a5246 = a5244 & ~i108;
assign a5248 = a5246 & i106;
assign a5250 = a5248 & l326;
assign a5252 = a5240 & ~a864;
assign a5254 = a5252 & ~i106;
assign a5256 = a5254 & ~i110;
assign a5258 = a5256 & i108;
assign a5260 = a5258 & l326;
assign a5262 = a3620 & ~l294;
assign a5264 = a5262 & l326;
assign a5266 = ~a5264 & ~a5260;
assign a5268 = a5266 & ~a5250;
assign a5270 = a5268 & ~a4388;
assign a5272 = a5270 & ~a5238;
assign a5274 = a5272 & ~a5110;
assign a5276 = a5274 & ~a3526;
assign a5278 = a5276 & ~a3638;
assign a5280 = a5278 & ~a3650;
assign a5282 = a5280 & ~a3662;
assign a5284 = a5282 & ~a3668;
assign a5286 = a5284 & ~a3674;
assign a5288 = a5286 & ~a3678;
assign a5290 = a5288 & ~a3680;
assign a5292 = a5290 & ~a3682;
assign a5294 = ~a5292 & a3710;
assign a5296 = a5294 & ~a5104;
assign a5298 = a5296 & ~a5090;
assign a5300 = a5298 & ~a5086;
assign a5302 = a5300 & ~a5078;
assign a5304 = a5302 & ~a5068;
assign a5306 = a3446 & ~a960;
assign a5308 = a5306 & i110;
assign a5310 = a5308 & ~i108;
assign a5312 = a5310 & ~i106;
assign a5314 = a3446 & ~l294;
assign a5316 = a5314 & ~a1062;
assign a5318 = a5316 & i110;
assign a5320 = a5318 & ~i108;
assign a5322 = a5320 & i106;
assign a5324 = a5314 & ~a864;
assign a5326 = a5324 & ~i106;
assign a5328 = a5326 & ~i110;
assign a5330 = a5328 & i108;
assign a5332 = a3724 & ~l294;
assign a5334 = ~a5332 & ~a5330;
assign a5336 = a5334 & ~a5322;
assign a5338 = a5336 & ~a5312;
assign a5340 = a5338 & ~a5304;
assign a5342 = a5340 & ~a5064;
assign a5344 = a5342 & ~a3454;
assign a5346 = a5052 & ~l284;
assign a5348 = a5346 & i112;
assign a5350 = a5348 & ~l236;
assign a5352 = a5054 & ~l286;
assign a5354 = a5352 & i114;
assign a5356 = ~a5354 & ~a5350;
assign a5358 = a5356 & ~a5344;
assign a5360 = a5358 & a3442;
assign a5362 = a5360 & ~a5058;
assign a5364 = ~a5362 & ~l274;
assign a5366 = ~a5364 & ~a2680;
assign a5368 = a5366 & ~a2678;
assign a5370 = a5368 & ~a2668;
assign a5372 = a5370 & ~a2656;
assign a5374 = a5372 & ~a2644;
assign a5376 = ~a5374 & ~a2640;
assign a5378 = a5376 & ~a2634;
assign a5380 = a5378 & ~a2626;
assign a5382 = a5380 & ~a2618;
assign a5384 = a5382 & ~a2616;
assign a5386 = a5384 & ~a2606;
assign a5388 = a5386 & ~a3416;
assign a5390 = a5388 & ~a2586;
assign a5392 = a5390 & ~a4330;
assign a5394 = a5392 & ~a2564;
assign a5396 = a5394 & ~a2550;
assign a5398 = a5396 & ~a2544;
assign a5400 = ~a5398 & ~a2538;
assign a5402 = ~a5400 & ~a2532;
assign a5404 = ~a5402 & ~a2516;
assign a5406 = a5404 & ~a2514;
assign a5408 = a5406 & ~a2504;
assign a5410 = a5408 & ~a2492;
assign a5412 = a5410 & ~a2488;
assign a5414 = ~a5412 & ~a2484;
assign a5416 = a5414 & ~a2478;
assign a5418 = a5416 & ~a2470;
assign a5420 = a5418 & ~a2462;
assign a5422 = a5420 & ~a2460;
assign a5424 = a5422 & ~a2458;
assign a5426 = a5424 & ~a3400;
assign a5428 = a5426 & ~a2438;
assign a5430 = a5428 & ~a4322;
assign a5432 = a5430 & ~a2416;
assign a5434 = a5432 & ~a2408;
assign a5436 = ~a5434 & ~a2402;
assign a5438 = a5436 & ~a2398;
assign a5440 = a5438 & ~a2392;
assign a5442 = a5440 & ~a2380;
assign a5444 = a5442 & ~a2378;
assign a5446 = ~a5444 & ~a2372;
assign a5448 = a5446 & ~a2368;
assign a5450 = a5448 & ~a2360;
assign a5452 = a5450 & ~a2352;
assign a5454 = a5452 & ~a2342;
assign a5456 = a5454 & ~a3392;
assign a5458 = a5456 & ~a2332;
assign a5460 = a5458 & ~a2324;
assign a5462 = a5460 & ~a2314;
assign a5464 = ~a5462 & ~a2302;
assign a5466 = a5464 & ~a2300;
assign a5468 = ~a5466 & ~a2294;
assign a5470 = a5468 & ~a2290;
assign a5472 = a5470 & ~a2282;
assign a5474 = a5472 & ~a2274;
assign a5476 = a5474 & ~a3386;
assign a5478 = a5476 & ~a2264;
assign a5480 = a5478 & ~a2256;
assign a5482 = ~a5480 & ~a2246;
assign a5484 = a5482 & ~a2234;
assign a5486 = ~a5484 & ~a2232;
assign a5488 = a5486 & ~a2226;
assign a5490 = a5488 & ~a2218;
assign a5492 = a5490 & ~a2210;
assign a5494 = a5492 & ~a2208;
assign a5496 = a5494 & ~a2206;
assign a5498 = ~a5496 & ~a2204;
assign a5500 = a5498 & ~a2198;
assign a5502 = ~a5500 & ~a2194;
assign a5504 = ~a5502 & ~a2188;
assign a5506 = a5504 & ~a2182;
assign a5508 = a5506 & ~a2168;
assign a5510 = a5508 & ~a2166;
assign a5512 = a5510 & ~a2164;
assign a5514 = a5512 & ~a2158;
assign a5516 = a5514 & ~a2156;
assign a5518 = a5516 & ~a2154;
assign a5520 = ~a5518 & ~a2146;
assign a5522 = a5520 & ~a2142;
assign a5524 = a5522 & ~a2134;
assign a5526 = a5524 & ~a2126;
assign a5528 = a5526 & ~a2124;
assign a5530 = ~a5528 & ~a2122;
assign a5532 = a5530 & ~a2118;
assign a5534 = a5532 & ~a2108;
assign a5536 = a5534 & ~a2096;
assign a5538 = a5536 & ~a2084;
assign a5540 = a5538 & ~a2076;
assign a5542 = a5540 & ~a2068;
assign a5544 = a5542 & ~a2054;
assign a5546 = a5544 & ~a2052;
assign a5548 = a5546 & ~a2042;
assign a5550 = a5548 & ~a2036;
assign a5552 = ~a5550 & ~a2032;
assign a5554 = a5552 & ~a2028;
assign a5556 = a5554 & ~a2020;
assign a5558 = a5556 & ~a2010;
assign a5560 = ~a5558 & ~a2008;
assign a5562 = a5560 & ~a2004;
assign a5564 = a5562 & ~a2000;
assign a5566 = a5564 & ~a1984;
assign a5568 = ~a5566 & ~a1980;
assign a5570 = a5568 & ~a1978;
assign a5572 = a5570 & ~a1976;
assign a5574 = a5572 & ~a1968;
assign a5576 = a5574 & ~a1966;
assign a5578 = ~a5576 & ~a1960;
assign a5580 = ~a5578 & ~a1950;
assign a5582 = a5580 & ~a1944;
assign a5584 = a5582 & ~a1938;
assign a5586 = a5584 & ~a1936;
assign a5588 = a5586 & ~a1934;
assign a5590 = a5588 & ~a1932;
assign a5592 = a5590 & ~a1930;
assign a5594 = ~a5592 & ~a1928;
assign a5596 = a5594 & ~a1916;
assign a5598 = a5596 & ~a1908;
assign a5600 = a5598 & ~a1892;
assign a5602 = ~a5600 & ~a1890;
assign a5604 = a5602 & ~a1884;
assign a5606 = a5604 & ~a1876;
assign a5608 = a5606 & ~a1866;
assign a5610 = a5608 & ~a3372;
assign a5612 = ~a5610 & ~a1850;
assign a5614 = ~a5612 & ~a1838;
assign a5616 = a5614 & ~a1834;
assign a5618 = a5616 & ~a1826;
assign a5620 = a5618 & ~a1824;
assign a5622 = a5620 & ~a3366;
assign a5624 = a5622 & ~a3364;
assign a5626 = a5624 & ~a3362;
assign a5628 = ~a5626 & ~a3360;
assign a5630 = a5628 & ~a1796;
assign a5632 = a5630 & ~a1786;
assign a5634 = a5632 & ~a1770;
assign a5636 = ~a5634 & ~a1768;
assign a5638 = a5636 & ~a1762;
assign a5640 = a5638 & ~a1754;
assign a5642 = a5640 & ~a1744;
assign a5644 = a5642 & ~a3354;
assign a5646 = ~a5644 & ~a1728;
assign a5648 = ~a5646 & ~a1716;
assign a5650 = a5648 & ~a1712;
assign a5652 = a5650 & ~a1704;
assign a5654 = a5652 & ~a1702;
assign a5656 = a5654 & ~a3348;
assign a5658 = a5656 & ~a3346;
assign a5660 = a5658 & ~a3344;
assign a5662 = ~a5660 & ~a3342;
assign a5664 = a5662 & ~a1674;
assign a5666 = a5664 & ~a1664;
assign a5668 = a5666 & ~a1648;
assign a5670 = ~a5668 & ~a1646;
assign a5672 = a5670 & ~a1640;
assign a5674 = a5672 & ~a1632;
assign a5676 = ~a5674 & ~a1624;
assign a5678 = ~a5676 & ~a1618;
assign a5680 = ~a5678 & ~a1606;
assign a5682 = ~a5680 & ~a1594;
assign a5684 = a5682 & ~a1590;
assign a5686 = a5684 & ~a1582;
assign a5688 = ~a5686 & ~a1574;
assign a5690 = a5688 & ~a1566;
assign a5692 = a5690 & ~a1558;
assign a5694 = a5692 & ~a1548;
assign a5696 = a5694 & ~a1538;
assign a5698 = a5696 & ~a1528;
assign a5700 = a5698 & ~a1522;
assign a5702 = ~a5700 & ~a1506;
assign a5704 = a5702 & ~a1502;
assign a5706 = a5704 & ~a1494;
assign a5708 = a5706 & ~a1486;
assign a5710 = a5708 & ~a1482;
assign a5712 = a5710 & ~a1478;
assign a5714 = a5712 & ~a1476;
assign a5716 = ~a5714 & ~a1472;
assign a5718 = a5716 & ~a1462;
assign a5720 = a5718 & ~a1448;
assign a5722 = a5720 & ~a1446;
assign a5724 = ~a5722 & ~a1442;
assign a5726 = a5724 & ~a1436;
assign a5728 = a5726 & ~a1428;
assign a5730 = a5728 & ~a1420;
assign a5732 = a5730 & ~a1418;
assign a5734 = a5732 & ~a1416;
assign a5736 = ~a5734 & ~a1414;
assign a5738 = a5736 & ~a1408;
assign a5740 = ~a5738 & ~a1404;
assign a5742 = ~a5740 & ~a1398;
assign a5744 = a5742 & ~a1392;
assign a5746 = a5744 & ~a1378;
assign a5748 = ~a5746 & ~a1376;
assign a5750 = a5748 & ~a1372;
assign a5752 = a5750 & ~a1364;
assign a5754 = a5752 & ~a1356;
assign a5756 = ~a5754 & ~a1352;
assign a5758 = a5756 & ~a1346;
assign a5760 = a5758 & ~a1338;
assign a5762 = a5760 & ~a1330;
assign a5764 = a5762 & ~a1320;
assign a5766 = a5764 & ~a1306;
assign a5768 = ~a5766 & ~a1290;
assign a5770 = a5768 & ~a1284;
assign a5772 = a5770 & ~a1278;
assign a5774 = a5772 & ~a1268;
assign a5776 = ~a5774 & ~a1254;
assign a5778 = a5776 & ~a1242;
assign a5780 = a5778 & ~a1230;
assign a5782 = a5780 & ~a1222;
assign a5784 = a5782 & ~a1214;
assign a5786 = a5784 & ~a1200;
assign a5788 = ~a5786 & ~a1198;
assign a5790 = a5788 & ~a1194;
assign a5792 = a5790 & ~a1186;
assign a5794 = a5792 & ~a1178;
assign a5796 = ~a5794 & ~a1176;
assign a5798 = ~a5796 & ~a4314;
assign a5800 = a5798 & ~a1162;
assign a5802 = a5800 & ~a1156;
assign a5804 = a5802 & ~a1152;
assign a5806 = a5804 & ~a1150;
assign a5808 = a5806 & ~a1140;
assign a5810 = a5808 & ~a1128;
assign a5812 = a5810 & ~a1116;
assign a5814 = ~a5812 & ~a1104;
assign a5816 = a5814 & ~a1100;
assign a5818 = a5816 & ~a1090;
assign a5820 = a5818 & ~a1080;
assign a5822 = ~a5820 & ~a1060;
assign a5824 = a5822 & ~a1056;
assign a5826 = a5824 & ~a1048;
assign a5828 = a5826 & ~a4306;
assign a5830 = a5828 & ~a1038;
assign a5832 = a5830 & ~a1032;
assign a5834 = ~a5832 & ~a1030;
assign a5836 = a5834 & ~a1024;
assign a5838 = a5836 & ~a1010;
assign a5840 = a5838 & ~a996;
assign a5842 = a5840 & ~a992;
assign a5844 = a5842 & ~a986;
assign a5846 = a5844 & ~a982;
assign a5848 = ~a5846 & ~a968;
assign a5850 = a5848 & ~a964;
assign a5852 = a5850 & ~a956;
assign a5854 = a5852 & ~a3322;
assign a5856 = a5854 & ~a3318;
assign a5858 = a5856 & ~a934;
assign a5860 = a5858 & ~a928;
assign a5862 = ~a5860 & ~a3314;
assign a5864 = ~a5862 & ~a4298;
assign a5866 = a5864 & ~a908;
assign a5868 = a5866 & ~a902;
assign a5870 = ~a5868 & ~a896;
assign a5872 = a5870 & ~a888;
assign a5874 = ~a5872 & ~a876;
assign a5876 = ~a5874 & ~a860;
assign a5878 = ~a5876 & i102;
assign a5880 = a5876 & ~i102;
assign a5882 = ~a5880 & ~a5878;
assign a5884 = a4294 & l304;
assign a5886 = a5884 & l326;
assign a5888 = a4304 & l302;
assign a5890 = a5888 & l304;
assign a5892 = a4348 & i64;
assign a5894 = a5892 & ~l294;
assign a5896 = a5894 & l326;
assign a5898 = a4348 & ~l294;
assign a5900 = a5898 & ~a864;
assign a5902 = a5900 & ~i110;
assign a5904 = a5902 & i108;
assign a5906 = a5904 & ~i106;
assign a5908 = a5906 & l326;
assign a5910 = a5898 & ~a1062;
assign a5912 = a5910 & i110;
assign a5914 = a5912 & ~i108;
assign a5916 = a5914 & i106;
assign a5918 = a5916 & l326;
assign a5920 = a5892 & a864;
assign a5922 = a5892 & a1062;
assign a5924 = a5892 & a1084;
assign a5926 = a5924 & ~l326;
assign a5928 = a4348 & a1062;
assign a5930 = a5928 & ~l330;
assign a5932 = a5930 & i156;
assign a5934 = a4348 & a864;
assign a5936 = a5934 & ~l330;
assign a5938 = a5936 & i156;
assign a5940 = a4348 & ~a1062;
assign a5942 = a5940 & i110;
assign a5944 = a5942 & ~i108;
assign a5946 = a5944 & i106;
assign a5948 = a5946 & ~l326;
assign a5950 = a5948 & l330;
assign a5952 = a4348 & ~a864;
assign a5954 = a5952 & ~i106;
assign a5956 = a5954 & ~i110;
assign a5958 = a5956 & i108;
assign a5960 = a5958 & ~l326;
assign a5962 = a5960 & l330;
assign a5964 = a4348 & l216;
assign a5966 = a5964 & ~i44;
assign a5968 = a4348 & ~a952;
assign a5970 = a5968 & i110;
assign a5972 = a5970 & i108;
assign a5974 = a5972 & ~i106;
assign a5976 = a4348 & ~a960;
assign a5978 = a5976 & i110;
assign a5980 = a5978 & ~i108;
assign a5982 = a5980 & ~i106;
assign a5984 = a4348 & ~l288;
assign a5986 = a5984 & l290;
assign a5988 = a5986 & ~i118;
assign a5990 = a5892 & l294;
assign a5992 = a5990 & l326;
assign a5994 = a4348 & l294;
assign a5996 = a5994 & ~a1062;
assign a5998 = a5996 & i110;
assign a6000 = a5998 & ~i108;
assign a6002 = a6000 & i106;
assign a6004 = a6002 & l326;
assign a6006 = a5994 & ~a864;
assign a6008 = a6006 & ~i106;
assign a6010 = a6008 & ~i110;
assign a6012 = a6010 & i108;
assign a6014 = a6012 & l326;
assign a6016 = a5984 & i116;
assign a6018 = a4380 & ~l238;
assign a6020 = a6018 & l290;
assign a6022 = a6020 & a1084;
assign a6024 = a6022 & ~l298;
assign a6026 = a6024 & i126;
assign a6028 = a1986 & ~l270;
assign a6030 = a6028 & ~l268;
assign a6032 = a4380 & l290;
assign a6034 = a6032 & a952;
assign a6036 = a6034 & ~l298;
assign a6038 = a6036 & i126;
assign a6040 = ~a5172 & ~a5166;
assign a6042 = a6040 & ~a5164;
assign a6044 = a4380 & i64;
assign a6046 = a6044 & l290;
assign a6048 = a6046 & a952;
assign a6050 = ~a6048 & ~a6042;
assign a6052 = a6050 & ~a6038;
assign a6054 = ~a6052 & ~a5182;
assign a6056 = a6054 & ~a5184;
assign a6058 = a6056 & ~a5186;
assign a6060 = a6058 & ~a5194;
assign a6062 = a6060 & ~a5200;
assign a6064 = a6062 & ~a5206;
assign a6066 = ~a6064 & a6030;
assign a6068 = a6066 & ~l236;
assign a6070 = a6068 & ~a6026;
assign a6072 = ~a6070 & ~l276;
assign a6074 = ~a6072 & ~a6016;
assign a6076 = ~a6074 & ~a6014;
assign a6078 = a6076 & ~a6004;
assign a6080 = a6078 & ~a5992;
assign a6082 = a6080 & ~a5988;
assign a6084 = a6082 & ~a5982;
assign a6086 = ~a6084 & ~a5974;
assign a6088 = ~a6086 & ~a5966;
assign a6090 = a6088 & ~a5962;
assign a6092 = a6090 & ~a5950;
assign a6094 = a6092 & ~a5938;
assign a6096 = a6094 & ~a5932;
assign a6098 = a6096 & ~a5926;
assign a6100 = a6098 & ~a5922;
assign a6102 = a6100 & ~a5920;
assign a6104 = ~a6102 & ~a5918;
assign a6106 = a6104 & ~a5908;
assign a6108 = a6106 & ~a5896;
assign a6110 = ~a6108 & ~a4354;
assign a6112 = ~a6110 & ~a2764;
assign a6114 = ~a6112 & ~a2762;
assign a6116 = a6114 & ~a4342;
assign a6118 = a6116 & ~a2744;
assign a6120 = a6118 & ~a2742;
assign a6122 = a6120 & ~a2736;
assign a6124 = ~a6122 & ~a2728;
assign a6126 = a6124 & ~a2720;
assign a6128 = a6126 & ~a2712;
assign a6130 = a6128 & ~a2702;
assign a6132 = ~a6130 & ~a2698;
assign a6134 = ~a6132 & ~a2694;
assign a6136 = ~a6134 & ~a2688;
assign a6138 = ~a6136 & ~a2680;
assign a6140 = ~a6138 & ~a2678;
assign a6142 = a6140 & ~a3424;
assign a6144 = a6142 & ~a2656;
assign a6146 = a6144 & ~a2644;
assign a6148 = a6146 & ~a2640;
assign a6150 = a6148 & ~a2634;
assign a6152 = ~a6150 & ~a2626;
assign a6154 = ~a6152 & ~a2618;
assign a6156 = a6154 & ~a2616;
assign a6158 = a6156 & ~a2606;
assign a6160 = a6158 & ~a3416;
assign a6162 = ~a6160 & ~a2586;
assign a6164 = a6162 & ~a2576;
assign a6166 = a6164 & ~a2564;
assign a6168 = a6166 & ~a2550;
assign a6170 = a6168 & ~a2544;
assign a6172 = a6170 & ~a2538;
assign a6174 = ~a6172 & ~a2532;
assign a6176 = ~a6174 & ~a2516;
assign a6178 = ~a6176 & ~a2514;
assign a6180 = a6178 & ~a3408;
assign a6182 = a6180 & ~a2492;
assign a6184 = a6182 & ~a2488;
assign a6186 = a6184 & ~a2484;
assign a6188 = a6186 & ~a2478;
assign a6190 = ~a6188 & ~a2470;
assign a6192 = ~a6190 & ~a2462;
assign a6194 = a6192 & ~a2460;
assign a6196 = a6194 & ~a2458;
assign a6198 = a6196 & ~a3400;
assign a6200 = ~a6198 & ~a2438;
assign a6202 = a6200 & ~a2428;
assign a6204 = a6202 & ~a2416;
assign a6206 = a6204 & ~a2408;
assign a6208 = ~a6206 & ~a2402;
assign a6210 = ~a6208 & ~a2398;
assign a6212 = ~a6210 & ~a2392;
assign a6214 = ~a6212 & ~a2380;
assign a6216 = ~a6214 & ~a2378;
assign a6218 = a6216 & ~a2372;
assign a6220 = a6218 & ~a2368;
assign a6222 = ~a6220 & ~a2360;
assign a6224 = ~a6222 & ~a2352;
assign a6226 = a6224 & ~a2342;
assign a6228 = a6226 & ~a3392;
assign a6230 = a6228 & ~a2332;
assign a6232 = ~a6230 & ~a2324;
assign a6234 = a6232 & ~a2314;
assign a6236 = a6234 & ~a2302;
assign a6238 = ~a6236 & ~a2300;
assign a6240 = a6238 & ~a2294;
assign a6242 = a6240 & ~a2290;
assign a6244 = ~a6242 & ~a2282;
assign a6246 = ~a6244 & ~a2274;
assign a6248 = a6246 & ~a3386;
assign a6250 = a6248 & ~a2264;
assign a6252 = ~a6250 & ~a2256;
assign a6254 = a6252 & ~a2246;
assign a6256 = a6254 & ~a2234;
assign a6258 = ~a6256 & ~a2232;
assign a6260 = a6258 & ~a2226;
assign a6262 = ~a6260 & ~a2218;
assign a6264 = ~a6262 & ~a2210;
assign a6266 = a6264 & ~a2208;
assign a6268 = a6266 & ~a2206;
assign a6270 = a6268 & ~a2204;
assign a6272 = a6270 & ~a2198;
assign a6274 = ~a6272 & ~a2194;
assign a6276 = a6274 & ~a2188;
assign a6278 = a6276 & ~a2182;
assign a6280 = a6278 & ~a2168;
assign a6282 = a6280 & ~a2166;
assign a6284 = a6282 & ~a2164;
assign a6286 = a6284 & ~a2158;
assign a6288 = a6286 & ~a2156;
assign a6290 = a6288 & ~a2154;
assign a6292 = ~a6290 & ~a2146;
assign a6294 = a6292 & ~a2142;
assign a6296 = ~a6294 & ~a2134;
assign a6298 = ~a6296 & ~a2126;
assign a6300 = a6298 & ~a2124;
assign a6302 = ~a6300 & ~a2122;
assign a6304 = a6302 & ~a2118;
assign a6306 = a6304 & ~a2108;
assign a6308 = a6306 & ~a2096;
assign a6310 = a6308 & ~a2084;
assign a6312 = a6310 & ~a2076;
assign a6314 = a6312 & ~a2068;
assign a6316 = ~a6314 & ~a2054;
assign a6318 = a6316 & ~a3380;
assign a6320 = a6318 & ~a2042;
assign a6322 = a6320 & ~a2036;
assign a6324 = a6322 & ~a2032;
assign a6326 = a6324 & ~a2028;
assign a6328 = ~a6326 & ~a2020;
assign a6330 = ~a6328 & ~a2010;
assign a6332 = ~a6330 & ~a2008;
assign a6334 = a6332 & ~a2004;
assign a6336 = a6334 & ~a2000;
assign a6338 = a6336 & ~a1984;
assign a6340 = ~a6338 & ~a1980;
assign a6342 = ~a6340 & ~a1978;
assign a6344 = ~a6342 & ~a1976;
assign a6346 = a6344 & ~a1968;
assign a6348 = a6346 & ~a1966;
assign a6350 = ~a6348 & ~a1960;
assign a6352 = ~a6350 & ~a1950;
assign a6354 = ~a6352 & ~a1944;
assign a6356 = ~a6354 & ~a1938;
assign a6358 = a6356 & ~a1936;
assign a6360 = a6358 & ~a1934;
assign a6362 = a6360 & ~a1932;
assign a6364 = a6362 & ~a1930;
assign a6366 = ~a6364 & ~a1928;
assign a6368 = a6366 & ~a1916;
assign a6370 = a6368 & ~a1908;
assign a6372 = a6370 & ~a1892;
assign a6374 = ~a6372 & ~a1890;
assign a6376 = ~a6374 & ~a1884;
assign a6378 = ~a6376 & ~a1876;
assign a6380 = a6378 & ~a1866;
assign a6382 = a6380 & ~a3372;
assign a6384 = ~a6382 & ~a1850;
assign a6386 = ~a6384 & ~a1838;
assign a6388 = ~a6386 & ~a1834;
assign a6390 = ~a6388 & ~a1826;
assign a6392 = a6390 & ~a1824;
assign a6394 = a6392 & ~a3366;
assign a6396 = a6394 & ~a3364;
assign a6398 = a6396 & ~a3362;
assign a6400 = ~a6398 & ~a3360;
assign a6402 = a6400 & ~a1796;
assign a6404 = a6402 & ~a1786;
assign a6406 = a6404 & ~a1770;
assign a6408 = ~a6406 & ~a1768;
assign a6410 = a6408 & ~a1762;
assign a6412 = a6410 & ~a1754;
assign a6414 = a6412 & ~a1744;
assign a6416 = a6414 & ~a3354;
assign a6418 = ~a6416 & ~a1728;
assign a6420 = ~a6418 & ~a1716;
assign a6422 = a6420 & ~a1712;
assign a6424 = a6422 & ~a1704;
assign a6426 = a6424 & ~a1702;
assign a6428 = a6426 & ~a3348;
assign a6430 = a6428 & ~a3346;
assign a6432 = a6430 & ~a3344;
assign a6434 = ~a6432 & ~a3342;
assign a6436 = a6434 & ~a1674;
assign a6438 = a6436 & ~a1664;
assign a6440 = a6438 & ~a1648;
assign a6442 = ~a6440 & ~a1646;
assign a6444 = a6442 & ~a1640;
assign a6446 = ~a6444 & ~a1632;
assign a6448 = ~a6446 & ~a1624;
assign a6450 = ~a6448 & ~a1618;
assign a6452 = a6450 & ~a1606;
assign a6454 = ~a6452 & ~a1594;
assign a6456 = a6454 & ~a1590;
assign a6458 = ~a6456 & ~a1582;
assign a6460 = a6458 & ~a1574;
assign a6462 = a6460 & ~a1566;
assign a6464 = a6462 & ~a1558;
assign a6466 = a6464 & ~a1548;
assign a6468 = a6466 & ~a1538;
assign a6470 = a6468 & ~a1528;
assign a6472 = a6470 & ~a1522;
assign a6474 = ~a6472 & ~a1506;
assign a6476 = a6474 & ~a1502;
assign a6478 = ~a6476 & ~a1494;
assign a6480 = ~a6478 & ~a1486;
assign a6482 = a6480 & ~a1482;
assign a6484 = a6482 & ~a1478;
assign a6486 = a6484 & ~a1476;
assign a6488 = ~a6486 & ~a1472;
assign a6490 = a6488 & ~a1462;
assign a6492 = a6490 & ~a1448;
assign a6494 = ~a6492 & ~a1446;
assign a6496 = a6494 & ~a1442;
assign a6498 = a6496 & ~a1436;
assign a6500 = ~a6498 & ~a1428;
assign a6502 = ~a6500 & ~a1420;
assign a6504 = a6502 & ~a1418;
assign a6506 = a6504 & ~a1416;
assign a6508 = a6506 & ~a1414;
assign a6510 = a6508 & ~a1408;
assign a6512 = ~a6510 & ~a1404;
assign a6514 = a6512 & ~a1398;
assign a6516 = a6514 & ~a1392;
assign a6518 = ~a6516 & ~a1378;
assign a6520 = a6518 & ~a1376;
assign a6522 = a6520 & ~a1372;
assign a6524 = ~a6522 & ~a1364;
assign a6526 = ~a6524 & ~a1356;
assign a6528 = a6526 & ~a1352;
assign a6530 = a6528 & ~a1346;
assign a6532 = a6530 & ~a1338;
assign a6534 = a6532 & ~a1330;
assign a6536 = a6534 & ~a1320;
assign a6538 = a6536 & ~a1306;
assign a6540 = ~a6538 & ~a1290;
assign a6542 = a6540 & ~a1284;
assign a6544 = a6542 & ~a1278;
assign a6546 = a6544 & ~a1268;
assign a6548 = a6546 & ~a1254;
assign a6550 = a6548 & ~a1242;
assign a6552 = a6550 & ~a1230;
assign a6554 = a6552 & ~a1222;
assign a6556 = a6554 & ~a1214;
assign a6558 = a6556 & ~a1200;
assign a6560 = ~a6558 & ~a1198;
assign a6562 = a6560 & ~a1194;
assign a6564 = ~a6562 & ~a1186;
assign a6566 = ~a6564 & ~a1178;
assign a6568 = ~a6566 & ~a1176;
assign a6570 = a6568 & ~a1172;
assign a6572 = a6570 & ~a1162;
assign a6574 = a6572 & ~a1156;
assign a6576 = a6574 & ~a1152;
assign a6578 = a6576 & ~a1150;
assign a6580 = a6578 & ~a1140;
assign a6582 = a6580 & ~a1128;
assign a6584 = a6582 & ~a1116;
assign a6586 = a6584 & ~a1104;
assign a6588 = a6586 & ~a1100;
assign a6590 = a6588 & ~a1090;
assign a6592 = a6590 & ~a1080;
assign a6594 = ~a6592 & ~a1060;
assign a6596 = a6594 & ~a1056;
assign a6598 = ~a6596 & ~a1048;
assign a6600 = a6598 & ~a1040;
assign a6602 = a6600 & ~a1038;
assign a6604 = a6602 & ~a1032;
assign a6606 = ~a6604 & ~a1030;
assign a6608 = a6606 & ~a5890;
assign a6610 = ~a6608 & ~a1010;
assign a6612 = ~a6610 & ~a3336;
assign a6614 = a6612 & ~a992;
assign a6616 = a6614 & ~a986;
assign a6618 = ~a6616 & ~a982;
assign a6620 = ~a6618 & ~a968;
assign a6622 = a6620 & ~a964;
assign a6624 = ~a6622 & ~a956;
assign a6626 = ~a6624 & ~a3322;
assign a6628 = a6626 & ~a3318;
assign a6630 = a6628 & ~a934;
assign a6632 = a6630 & ~a928;
assign a6634 = ~a6632 & ~a3314;
assign a6636 = a6634 & ~a912;
assign a6638 = a6636 & ~a908;
assign a6640 = a6638 & ~a902;
assign a6642 = ~a6640 & ~a5886;
assign a6644 = a6642 & ~a888;
assign a6646 = ~a6644 & ~a876;
assign a6648 = a6646 & ~a860;
assign a6650 = ~a6648 & i104;
assign a6652 = a6648 & ~i104;
assign a6654 = ~a6652 & ~a6650;
assign a6656 = l258 & ~l256;
assign a6658 = a6656 & ~l254;
assign a6660 = ~l252 & l250;
assign a6662 = a6660 & l248;
assign a6664 = a6662 & l236;
assign a6666 = a6664 & ~l184;
assign a6668 = a6666 & l260;
assign a6670 = a6668 & l262;
assign a6672 = a6670 & a6658;
assign a6674 = a6672 & ~l240;
assign a6676 = l246 & ~l244;
assign a6678 = a6676 & l242;
assign a6680 = a6678 & a6674;
assign a6682 = a6680 & ~l266;
assign a6684 = a6682 & i94;
assign a6686 = l258 & l256;
assign a6688 = a6686 & ~l254;
assign a6690 = a6688 & a6670;
assign a6692 = a6690 & ~l240;
assign a6694 = a6692 & a6678;
assign a6696 = a6694 & ~l266;
assign a6698 = a6696 & i94;
assign a6700 = a6662 & ~l236;
assign a6702 = a6700 & ~l238;
assign a6704 = a6702 & ~l184;
assign a6706 = a6704 & l260;
assign a6708 = a6706 & l262;
assign a6710 = a6708 & a6688;
assign a6712 = a6710 & ~l240;
assign a6714 = a6712 & a6678;
assign a6716 = a6714 & ~l266;
assign a6718 = a6716 & i94;
assign a6720 = l172 & l170;
assign a6722 = a6720 & ~l168;
assign a6724 = a6722 & ~l166;
assign a6726 = a6724 & ~l164;
assign a6728 = ~l258 & ~l256;
assign a6730 = a6728 & ~l254;
assign a6732 = a6664 & l260;
assign a6734 = a6732 & l262;
assign a6736 = a6734 & a6730;
assign a6738 = a6736 & ~l266;
assign a6740 = a6738 & i94;
assign a6742 = a6740 & a6726;
assign a6744 = a6662 & l184;
assign a6746 = a6744 & ~i12;
assign a6748 = a6746 & l260;
assign a6750 = a6748 & l262;
assign a6752 = a6750 & a6730;
assign a6754 = a6752 & ~l240;
assign a6756 = a6754 & ~l234;
assign a6758 = a6662 & ~l184;
assign a6760 = a6758 & ~l260;
assign a6762 = a6760 & i88;
assign a6764 = a6762 & l262;
assign a6766 = a6764 & a6730;
assign a6768 = a6766 & ~l240;
assign a6770 = a6768 & ~l234;
assign a6772 = a6758 & l260;
assign a6774 = a6772 & ~l262;
assign a6776 = a6774 & i90;
assign a6778 = a6776 & a6730;
assign a6780 = a6778 & ~l240;
assign a6782 = a6780 & ~l234;
assign a6784 = a6772 & l262;
assign a6786 = a6784 & ~a6730;
assign a6788 = a6786 & ~i86;
assign a6790 = a6788 & ~i84;
assign a6792 = a6790 & ~i82;
assign a6794 = a6792 & ~l240;
assign a6796 = a6794 & ~l234;
assign a6798 = a6784 & a6730;
assign a6800 = a6798 & l240;
assign a6802 = a6800 & ~i68;
assign a6804 = a6802 & ~l234;
assign a6806 = a6798 & ~l240;
assign a6808 = a6806 & l234;
assign a6810 = a6808 & ~i62;
assign a6812 = a6728 & l254;
assign a6814 = a6812 & a6670;
assign a6816 = a6814 & ~l240;
assign a6818 = a6816 & ~l266;
assign a6820 = a6818 & i94;
assign a6822 = a6820 & ~l234;
assign a6824 = a6664 & l184;
assign a6826 = a6824 & l260;
assign a6828 = a6826 & l262;
assign a6830 = a6828 & a6812;
assign a6832 = a6830 & ~l240;
assign a6834 = ~l246 & l244;
assign a6836 = a6834 & l242;
assign a6838 = a6836 & a6832;
assign a6840 = a6838 & ~l266;
assign a6842 = a6840 & i94;
assign a6844 = a6842 & ~l234;
assign a6846 = a6660 & ~l248;
assign a6848 = a6846 & l236;
assign a6850 = a6848 & ~i64;
assign a6852 = a6846 & ~l234;
assign a6854 = a6852 & i62;
assign a6856 = a6846 & ~a6836;
assign a6858 = ~i74 & i70;
assign a6860 = a6858 & i72;
assign a6862 = a6860 & a6856;
assign a6864 = a6846 & ~l240;
assign a6866 = a6864 & i68;
assign a6868 = a6846 & ~l184;
assign a6870 = a6868 & i12;
assign a6872 = a6846 & l260;
assign a6874 = a6872 & ~i88;
assign a6876 = a6846 & l262;
assign a6878 = a6876 & ~i90;
assign a6880 = a6846 & ~a6688;
assign a6882 = i86 & i84;
assign a6884 = a6882 & ~i82;
assign a6886 = a6884 & a6880;
assign a6888 = a6846 & ~a6812;
assign a6890 = ~i86 & i82;
assign a6892 = a6890 & ~i84;
assign a6894 = a6892 & a6888;
assign a6896 = ~l258 & l256;
assign a6898 = a6896 & ~l254;
assign a6900 = ~a6898 & a6846;
assign a6902 = ~i86 & i84;
assign a6904 = a6902 & ~i82;
assign a6906 = a6904 & a6900;
assign a6908 = a6846 & ~l264;
assign a6910 = a6908 & i92;
assign a6912 = a6846 & ~l266;
assign a6914 = a6912 & i94;
assign a6916 = a6846 & ~l232;
assign a6918 = a6916 & i60;
assign a6920 = a6846 & ~a6730;
assign a6922 = a6920 & ~i86;
assign a6924 = a6922 & ~i84;
assign a6926 = a6924 & ~i82;
assign a6928 = ~l252 & ~l250;
assign a6930 = a6928 & l248;
assign a6932 = a6930 & l236;
assign a6934 = a6932 & ~i64;
assign a6936 = a6934 & l238;
assign a6938 = a6930 & ~l236;
assign a6940 = a6938 & l238;
assign a6942 = a6940 & ~i66;
assign a6944 = a6930 & ~l234;
assign a6946 = a6944 & i62;
assign a6948 = a6930 & ~a6836;
assign a6950 = a6948 & i70;
assign a6952 = a6950 & ~i74;
assign a6954 = a6952 & i72;
assign a6956 = a6930 & ~l240;
assign a6958 = a6956 & i68;
assign a6960 = a6930 & ~l184;
assign a6962 = a6960 & i12;
assign a6964 = a6930 & l260;
assign a6966 = a6964 & ~i88;
assign a6968 = a6930 & l262;
assign a6970 = a6968 & ~i90;
assign a6972 = a6930 & ~a6658;
assign a6974 = i86 & ~i84;
assign a6976 = a6974 & ~i82;
assign a6978 = a6976 & a6972;
assign a6980 = a6930 & ~a6812;
assign a6982 = a6980 & i82;
assign a6984 = a6982 & ~i86;
assign a6986 = a6984 & ~i84;
assign a6988 = a6930 & ~a6898;
assign a6990 = a6988 & ~i86;
assign a6992 = a6990 & i84;
assign a6994 = a6992 & ~i82;
assign a6996 = a6930 & ~l264;
assign a6998 = a6996 & i92;
assign a7000 = a6930 & ~l266;
assign a7002 = a7000 & i94;
assign a7004 = a6930 & ~l232;
assign a7006 = a7004 & i60;
assign a7008 = a6930 & ~a6730;
assign a7010 = a7008 & ~i86;
assign a7012 = a7010 & ~i84;
assign a7014 = a7012 & ~i82;
assign a7016 = l252 & ~l250;
assign a7018 = a7016 & ~l248;
assign a7020 = a7018 & ~l234;
assign a7022 = a7020 & i62;
assign a7024 = a7018 & ~l240;
assign a7026 = a7024 & i68;
assign a7028 = a7018 & ~l184;
assign a7030 = a7028 & i12;
assign a7032 = a7018 & l260;
assign a7034 = a7032 & ~i88;
assign a7036 = a7018 & l262;
assign a7038 = a7036 & ~i90;
assign a7040 = a7018 & a6730;
assign a7042 = ~i86 & ~i84;
assign a7044 = a7042 & ~i82;
assign a7046 = ~a7044 & a7040;
assign a7048 = a7018 & ~l264;
assign a7050 = a7048 & i92;
assign a7052 = a7018 & ~l266;
assign a7054 = a7052 & i94;
assign a7056 = a7018 & ~l232;
assign a7058 = a7056 & i60;
assign a7060 = a6928 & ~l248;
assign a7062 = a7060 & l236;
assign a7064 = a7062 & ~i64;
assign a7066 = a7060 & a6726;
assign a7068 = i10 & i8;
assign a7070 = a7068 & ~i6;
assign a7072 = a7070 & ~i4;
assign a7074 = a7072 & ~i2;
assign a7076 = ~a7074 & a7066;
assign a7078 = a7060 & ~l240;
assign a7080 = a7078 & i68;
assign a7082 = a7060 & ~l184;
assign a7084 = a7082 & i12;
assign a7086 = a7060 & l260;
assign a7088 = a7086 & ~i88;
assign a7090 = a7060 & l262;
assign a7092 = a7090 & ~i90;
assign a7094 = a7060 & a6730;
assign a7096 = a7094 & ~a7044;
assign a7098 = a7060 & ~l264;
assign a7100 = a7098 & i92;
assign a7102 = a7060 & ~l232;
assign a7104 = a7102 & i60;
assign a7106 = l252 & l250;
assign a7108 = a7106 & ~l248;
assign a7110 = a7108 & ~l234;
assign a7112 = a7110 & i62;
assign a7114 = a7108 & ~l240;
assign a7116 = a7114 & i68;
assign a7118 = a7108 & ~l184;
assign a7120 = a7118 & i12;
assign a7122 = a7108 & l260;
assign a7124 = a7122 & ~i88;
assign a7126 = a7108 & l262;
assign a7128 = a7126 & ~i90;
assign a7130 = a7108 & a6730;
assign a7132 = a7130 & ~a7044;
assign a7134 = a7108 & ~l266;
assign a7136 = a7134 & i94;
assign a7138 = a7108 & ~l232;
assign a7140 = a7138 & i60;
assign a7142 = a7108 & ~l264;
assign a7144 = a7142 & i92;
assign a7146 = a7016 & l248;
assign a7148 = a7146 & ~a6730;
assign a7150 = a7016 & ~l264;
assign a7152 = a7150 & i92;
assign a7154 = a7016 & ~a6898;
assign a7156 = a7154 & ~i86;
assign a7158 = a7156 & i84;
assign a7160 = a7158 & ~i82;
assign a7162 = a7016 & ~a6688;
assign a7164 = a7162 & i86;
assign a7166 = a7164 & i84;
assign a7168 = a7166 & ~i82;
assign a7170 = a7016 & ~a6658;
assign a7172 = a7170 & i86;
assign a7174 = a7172 & ~i84;
assign a7176 = a7174 & ~i82;
assign a7178 = a7016 & l262;
assign a7180 = a7178 & ~i90;
assign a7182 = a7016 & l260;
assign a7184 = a7182 & ~i88;
assign a7186 = a7016 & ~l184;
assign a7188 = a7186 & i12;
assign a7190 = a7016 & ~l240;
assign a7192 = a7190 & i68;
assign a7194 = a7016 & ~l234;
assign a7196 = a7194 & i62;
assign a7198 = ~a7196 & ~a7192;
assign a7200 = a7198 & ~a7188;
assign a7202 = a7200 & ~a7184;
assign a7204 = a7202 & ~a7180;
assign a7206 = a7204 & ~a7176;
assign a7208 = a7206 & ~a7168;
assign a7210 = a7208 & ~a7160;
assign a7212 = a7210 & ~a7152;
assign a7214 = a7212 & a7148;
assign a7216 = a7214 & ~i86;
assign a7218 = a7216 & ~i84;
assign a7220 = a7218 & ~i82;
assign a7222 = ~a7220 & l248;
assign a7224 = a7222 & ~a7144;
assign a7226 = a7224 & ~a7140;
assign a7228 = a7226 & ~a7136;
assign a7230 = ~a7228 & ~a7132;
assign a7232 = a7230 & ~a7128;
assign a7234 = a7232 & ~a7124;
assign a7236 = a7234 & ~a7120;
assign a7238 = a7236 & ~a7116;
assign a7240 = a7238 & ~a7112;
assign a7242 = a7240 & ~a7104;
assign a7244 = a7242 & ~a7100;
assign a7246 = a7244 & ~a7096;
assign a7248 = a7246 & ~a7092;
assign a7250 = a7248 & ~a7088;
assign a7252 = a7250 & ~a7084;
assign a7254 = a7252 & ~a7080;
assign a7256 = a7254 & ~a7076;
assign a7258 = a7256 & ~a7064;
assign a7260 = ~a7258 & ~a7058;
assign a7262 = a7260 & ~a7054;
assign a7264 = ~a7262 & ~a7050;
assign a7266 = a7264 & ~a7046;
assign a7268 = a7266 & ~a7038;
assign a7270 = a7268 & ~a7034;
assign a7272 = a7270 & ~a7030;
assign a7274 = a7272 & ~a7026;
assign a7276 = a7274 & ~a7022;
assign a7278 = ~a7276 & ~a7014;
assign a7280 = ~a7278 & ~a7006;
assign a7282 = a7280 & ~a7002;
assign a7284 = a7282 & ~a6998;
assign a7286 = a7284 & ~a6994;
assign a7288 = a7286 & ~a6986;
assign a7290 = a7288 & ~a6978;
assign a7292 = a7290 & ~a6970;
assign a7294 = a7292 & ~a6966;
assign a7296 = a7294 & ~a6962;
assign a7298 = a7296 & ~a6958;
assign a7300 = a7298 & ~a6954;
assign a7302 = a7300 & ~a6946;
assign a7304 = a7302 & ~a6942;
assign a7306 = a7304 & ~a6936;
assign a7308 = ~a7306 & ~a6926;
assign a7310 = a7308 & ~a6918;
assign a7312 = a7310 & ~a6914;
assign a7314 = ~a7312 & ~a6910;
assign a7316 = a7314 & ~a6906;
assign a7318 = a7316 & ~a6894;
assign a7320 = a7318 & ~a6886;
assign a7322 = a7320 & ~a6878;
assign a7324 = a7322 & ~a6874;
assign a7326 = a7324 & ~a6870;
assign a7328 = a7326 & ~a6866;
assign a7330 = a7328 & ~a6862;
assign a7332 = a7330 & ~a6854;
assign a7334 = a7332 & ~a6850;
assign a7336 = a7334 & ~a6844;
assign a7338 = a7336 & ~a6822;
assign a7340 = ~a7338 & ~a6810;
assign a7342 = a7340 & ~a6804;
assign a7344 = a7342 & ~a6796;
assign a7346 = a7344 & ~a6782;
assign a7348 = a7346 & ~a6770;
assign a7350 = a7348 & ~a6756;
assign a7352 = a7350 & ~a6742;
assign a7354 = ~a7352 & ~a6718;
assign a7356 = a7354 & ~a6698;
assign a7358 = ~a7356 & ~a6684;
assign a7360 = ~a7358 & i76;
assign a7362 = a7358 & ~i76;
assign a7364 = ~a7362 & ~a7360;
assign a7366 = ~i86 & ~i82;
assign a7368 = a7366 & ~i84;
assign a7370 = a7368 & a6786;
assign a7372 = a7370 & ~l240;
assign a7374 = a7372 & ~l234;
assign a7376 = a6920 & ~i82;
assign a7378 = a7376 & ~i86;
assign a7380 = a7378 & ~i84;
assign a7382 = a7008 & ~i82;
assign a7384 = a7382 & ~i86;
assign a7386 = a7384 & ~i84;
assign a7388 = a7146 & ~l234;
assign a7390 = a7388 & i62;
assign a7392 = a7146 & ~l240;
assign a7394 = a7392 & i68;
assign a7396 = a7146 & ~l184;
assign a7398 = a7396 & i12;
assign a7400 = a7146 & l260;
assign a7402 = a7400 & ~i88;
assign a7404 = a7146 & l262;
assign a7406 = a7404 & ~i90;
assign a7408 = a7146 & ~a6658;
assign a7410 = a7408 & i86;
assign a7412 = a7410 & ~i84;
assign a7414 = a7412 & ~i82;
assign a7416 = a7146 & ~a6688;
assign a7418 = a7416 & i86;
assign a7420 = a7418 & i84;
assign a7422 = a7420 & ~i82;
assign a7424 = a7146 & ~a6898;
assign a7426 = a7424 & ~i86;
assign a7428 = a7426 & i84;
assign a7430 = a7428 & ~i82;
assign a7432 = a7146 & ~l264;
assign a7434 = a7432 & i92;
assign a7436 = a7148 & ~i82;
assign a7438 = a7436 & ~i86;
assign a7440 = a7438 & ~i84;
assign a7442 = ~a7440 & ~l250;
assign a7444 = a7442 & ~a7434;
assign a7446 = a7444 & ~a7430;
assign a7448 = a7446 & ~a7422;
assign a7450 = a7448 & ~a7414;
assign a7452 = a7450 & ~a7406;
assign a7454 = a7452 & ~a7402;
assign a7456 = a7454 & ~a7398;
assign a7458 = a7456 & ~a7394;
assign a7460 = a7458 & ~a7390;
assign a7462 = a7460 & ~a7144;
assign a7464 = a7462 & ~a7140;
assign a7466 = ~a7464 & ~a7136;
assign a7468 = ~a7466 & ~a7132;
assign a7470 = a7468 & ~a7128;
assign a7472 = a7470 & ~a7124;
assign a7474 = a7472 & ~a7120;
assign a7476 = a7474 & ~a7116;
assign a7478 = a7476 & ~a7112;
assign a7480 = a7478 & ~a7104;
assign a7482 = a7480 & ~a7100;
assign a7484 = a7482 & ~a7096;
assign a7486 = a7484 & ~a7092;
assign a7488 = a7486 & ~a7088;
assign a7490 = a7488 & ~a7084;
assign a7492 = a7490 & ~a7080;
assign a7494 = a7492 & ~a7076;
assign a7496 = a7494 & ~a7064;
assign a7498 = a7496 & ~a7058;
assign a7500 = a7498 & ~a7054;
assign a7502 = a7500 & ~a7050;
assign a7504 = a7502 & ~a7046;
assign a7506 = a7504 & ~a7038;
assign a7508 = a7506 & ~a7034;
assign a7510 = a7508 & ~a7030;
assign a7512 = a7510 & ~a7026;
assign a7514 = a7512 & ~a7022;
assign a7516 = a7514 & ~a7386;
assign a7518 = ~a7516 & ~a7006;
assign a7520 = a7518 & ~a7002;
assign a7522 = ~a7520 & ~a6998;
assign a7524 = a7522 & ~a6994;
assign a7526 = a7524 & ~a6986;
assign a7528 = a7526 & ~a6978;
assign a7530 = a7528 & ~a6970;
assign a7532 = a7530 & ~a6966;
assign a7534 = a7532 & ~a6962;
assign a7536 = a7534 & ~a6958;
assign a7538 = a7536 & ~a6954;
assign a7540 = a7538 & ~a6946;
assign a7542 = a7540 & ~a6942;
assign a7544 = a7542 & ~a6936;
assign a7546 = a7544 & ~a7380;
assign a7548 = a7546 & ~a6918;
assign a7550 = a7548 & ~a6914;
assign a7552 = a7550 & ~a6910;
assign a7554 = a7552 & ~a6906;
assign a7556 = a7554 & ~a6894;
assign a7558 = a7556 & ~a6886;
assign a7560 = a7558 & ~a6878;
assign a7562 = a7560 & ~a6874;
assign a7564 = a7562 & ~a6870;
assign a7566 = a7564 & ~a6866;
assign a7568 = a7566 & ~a6862;
assign a7570 = a7568 & ~a6854;
assign a7572 = a7570 & ~a6850;
assign a7574 = ~a7572 & ~a6844;
assign a7576 = a7574 & ~a6822;
assign a7578 = ~a7576 & ~a6810;
assign a7580 = a7578 & ~a6804;
assign a7582 = a7580 & ~a7374;
assign a7584 = a7582 & ~a6782;
assign a7586 = a7584 & ~a6770;
assign a7588 = a7586 & ~a6756;
assign a7590 = ~a7588 & ~a6742;
assign a7592 = a7590 & ~a6718;
assign a7594 = a7592 & ~a6698;
assign a7596 = ~a7594 & ~a6684;
assign a7598 = a7596 & i78;
assign a7600 = ~a7596 & ~i78;
assign a7602 = ~a7600 & ~a7598;
assign a7604 = ~i74 & i72;
assign a7606 = a7604 & i70;
assign a7608 = a7606 & a6856;
assign a7610 = a7042 & i82;
assign a7612 = a7610 & a6888;
assign a7614 = a6948 & ~i74;
assign a7616 = a7614 & i72;
assign a7618 = a7616 & i70;
assign a7620 = a6980 & ~i86;
assign a7622 = a7620 & ~i84;
assign a7624 = a7622 & i82;
assign a7626 = ~l250 & ~l248;
assign a7628 = a7626 & ~l232;
assign a7630 = a7628 & i60;
assign a7632 = l250 & ~l248;
assign a7634 = a7632 & a6730;
assign a7636 = a7634 & ~a7044;
assign a7638 = a7632 & ~l266;
assign a7640 = a7638 & i94;
assign a7642 = a7632 & ~l232;
assign a7644 = a7642 & i60;
assign a7646 = a7632 & ~l264;
assign a7648 = a7646 & i92;
assign a7650 = a6904 & ~a6898;
assign a7652 = ~l264 & i92;
assign a7654 = a6884 & ~a6688;
assign a7656 = a6976 & ~a6658;
assign a7658 = l262 & ~i90;
assign a7660 = l260 & ~i88;
assign a7662 = ~l184 & i12;
assign a7664 = ~l240 & i68;
assign a7666 = ~l234 & i62;
assign a7668 = ~a7666 & ~a7664;
assign a7670 = a7668 & ~a7662;
assign a7672 = a7670 & ~a7660;
assign a7674 = a7672 & ~a7658;
assign a7676 = a7674 & ~a7656;
assign a7678 = a7676 & ~a7654;
assign a7680 = a7678 & ~a7652;
assign a7682 = a7680 & ~a7650;
assign a7684 = ~l250 & l248;
assign a7686 = a7684 & ~a7682;
assign a7688 = a7686 & ~a7648;
assign a7690 = a7688 & ~a7644;
assign a7692 = a7690 & ~a7640;
assign a7694 = a7632 & l262;
assign a7696 = a7694 & ~i90;
assign a7698 = a7632 & l260;
assign a7700 = a7698 & ~i88;
assign a7702 = a7632 & ~l184;
assign a7704 = a7702 & i12;
assign a7706 = a7632 & ~l240;
assign a7708 = a7706 & i68;
assign a7710 = a7632 & ~l234;
assign a7712 = a7710 & i62;
assign a7714 = ~a7712 & ~a7708;
assign a7716 = a7714 & ~a7704;
assign a7718 = a7716 & ~a7700;
assign a7720 = a7718 & ~a7696;
assign a7722 = a7720 & ~a7692;
assign a7724 = a7722 & ~a7636;
assign a7726 = ~a7724 & l252;
assign a7728 = ~a7726 & ~a7104;
assign a7730 = a7728 & ~a7100;
assign a7732 = a7730 & ~a7096;
assign a7734 = a7732 & ~a7092;
assign a7736 = a7734 & ~a7088;
assign a7738 = a7736 & ~a7084;
assign a7740 = a7738 & ~a7080;
assign a7742 = a7740 & ~a7076;
assign a7744 = a7742 & ~a7064;
assign a7746 = a7626 & ~l266;
assign a7748 = a7746 & i94;
assign a7750 = ~a7748 & ~a7744;
assign a7752 = a7750 & ~a7630;
assign a7754 = ~a7752 & l252;
assign a7756 = a7754 & ~a7050;
assign a7758 = a7756 & ~a7046;
assign a7760 = a7758 & ~a7038;
assign a7762 = a7760 & ~a7034;
assign a7764 = a7762 & ~a7030;
assign a7766 = a7764 & ~a7026;
assign a7768 = a7766 & ~a7022;
assign a7770 = ~a7768 & ~a7386;
assign a7772 = ~a7770 & ~a7006;
assign a7774 = a7772 & ~a7002;
assign a7776 = a7774 & ~a6998;
assign a7778 = a7776 & ~a6994;
assign a7780 = a7778 & ~a7624;
assign a7782 = a7780 & ~a6978;
assign a7784 = a7782 & ~a6970;
assign a7786 = a7784 & ~a6966;
assign a7788 = a7786 & ~a6962;
assign a7790 = a7788 & ~a6958;
assign a7792 = a7790 & ~a7618;
assign a7794 = a7792 & ~a6946;
assign a7796 = a7794 & ~a6942;
assign a7798 = a7796 & ~a6936;
assign a7800 = ~a7798 & ~a7380;
assign a7802 = ~a7800 & ~a6918;
assign a7804 = a7802 & ~a6914;
assign a7806 = a7804 & ~a6910;
assign a7808 = a7806 & ~a6906;
assign a7810 = a7808 & ~a7612;
assign a7812 = a7810 & ~a6886;
assign a7814 = a7812 & ~a6878;
assign a7816 = a7814 & ~a6874;
assign a7818 = a7816 & ~a6870;
assign a7820 = a7818 & ~a6866;
assign a7822 = a7820 & ~a7608;
assign a7824 = a7822 & ~a6854;
assign a7826 = a7824 & ~a6850;
assign a7828 = ~a7826 & ~a6844;
assign a7830 = a7828 & ~a6822;
assign a7832 = a7830 & ~a6810;
assign a7834 = a7832 & ~a6804;
assign a7836 = a7834 & ~a7374;
assign a7838 = a7836 & ~a6782;
assign a7840 = a7838 & ~a6770;
assign a7842 = a7840 & ~a6756;
assign a7844 = ~a7842 & ~a6742;
assign a7846 = a7844 & ~a6718;
assign a7848 = a7846 & ~a6698;
assign a7850 = a7848 & ~a6684;
assign a7852 = ~a7850 & i80;
assign a7854 = a7850 & ~i80;
assign a7856 = ~a7854 & ~a7852;
assign a7858 = ~l172 & ~l170;
assign a7860 = a7858 & l168;
assign a7862 = a7860 & ~l166;
assign a7864 = a7862 & l164;
assign a7866 = a7864 & ~l236;
assign a7868 = a7866 & i64;
assign a7870 = a7868 & ~l234;
assign a7872 = a7864 & l236;
assign a7874 = a7872 & l240;
assign a7876 = a7874 & ~i68;
assign a7878 = a7876 & ~l234;
assign a7880 = a7872 & l234;
assign a7882 = a7880 & ~i62;
assign a7884 = a7872 & ~l198;
assign a7886 = a7884 & i26;
assign a7888 = a7886 & ~l234;
assign a7890 = a7872 & ~l200;
assign a7892 = a7890 & i28;
assign a7894 = a7892 & ~l234;
assign a7896 = a7872 & ~l202;
assign a7898 = a7896 & i30;
assign a7900 = a7898 & ~l234;
assign a7902 = a7872 & ~l204;
assign a7904 = a7902 & i32;
assign a7906 = a7904 & ~l234;
assign a7908 = a7872 & ~l206;
assign a7910 = a7908 & i34;
assign a7912 = a7910 & ~l234;
assign a7914 = a7872 & ~l196;
assign a7916 = a7914 & i24;
assign a7918 = a7916 & ~l234;
assign a7920 = a7868 & l234;
assign a7922 = ~l246 & ~l244;
assign a7924 = a7922 & ~l242;
assign a7926 = ~a7924 & a7872;
assign a7928 = a356 & ~i70;
assign a7930 = a7928 & a7926;
assign a7932 = a6676 & ~l242;
assign a7934 = ~a7932 & a7872;
assign a7936 = a7934 & a354;
assign a7938 = a6834 & ~l242;
assign a7940 = ~a7938 & a7872;
assign a7942 = ~i74 & ~i70;
assign a7944 = a7942 & i72;
assign a7946 = a7944 & a7940;
assign a7948 = l246 & l244;
assign a7950 = a7948 & ~l242;
assign a7952 = ~a7950 & a7872;
assign a7954 = i74 & i72;
assign a7956 = a7954 & ~i70;
assign a7958 = a7956 & a7952;
assign a7960 = a7922 & l242;
assign a7962 = ~a7960 & a7872;
assign a7964 = a7962 & a358;
assign a7966 = a7872 & l186;
assign a7968 = a7966 & ~i14;
assign a7970 = a7968 & l234;
assign a7972 = a7892 & l234;
assign a7974 = a7910 & l234;
assign a7976 = a7916 & l234;
assign a7978 = a7872 & ~l210;
assign a7980 = a7978 & i38;
assign a7982 = a7980 & l214;
assign a7984 = a7982 & ~l228;
assign a7986 = a7984 & l234;
assign a7988 = a7872 & l210;
assign a7990 = a7988 & ~l214;
assign a7992 = a7990 & i42;
assign a7994 = a7992 & ~l228;
assign a7996 = a7994 & l234;
assign a7998 = a7864 & ~l208;
assign a8000 = a7998 & i36;
assign a8002 = a8000 & l198;
assign a8004 = l172 & ~l170;
assign a8006 = a8004 & l168;
assign a8008 = a8006 & l166;
assign a8010 = a8008 & ~l164;
assign a8012 = a8010 & l240;
assign a8014 = a8012 & l198;
assign a8016 = l182 & ~l180;
assign a8018 = a8016 & l178;
assign a8020 = a8018 & l176;
assign a8022 = a8020 & ~l174;
assign a8024 = ~a8022 & a8014;
assign a8026 = a8024 & a8010;
assign a8028 = a8010 & ~l240;
assign a8030 = a8028 & l198;
assign a8032 = a8030 & ~a8022;
assign a8034 = a8032 & a8010;
assign a8036 = a8028 & ~l186;
assign a8038 = a8036 & ~a8022;
assign a8040 = a8038 & l172;
assign a8042 = a8040 & ~l170;
assign a8044 = a8042 & l168;
assign a8046 = a8044 & l166;
assign a8048 = a8046 & ~l164;
assign a8050 = a8012 & l186;
assign a8052 = a8050 & ~l198;
assign a8054 = a8052 & ~a8022;
assign a8056 = a8054 & l172;
assign a8058 = a8056 & ~l170;
assign a8060 = a8058 & l168;
assign a8062 = a8060 & l166;
assign a8064 = a8062 & ~l164;
assign a8066 = a8028 & l186;
assign a8068 = a8066 & ~l198;
assign a8070 = a8068 & ~a8022;
assign a8072 = a8070 & l172;
assign a8074 = a8072 & ~l170;
assign a8076 = a8074 & l168;
assign a8078 = a8076 & l166;
assign a8080 = a8078 & ~l164;
assign a8082 = a6724 & l164;
assign a8084 = a8082 & ~l214;
assign a8086 = a8084 & a7932;
assign a8088 = l182 & l180;
assign a8090 = a8088 & ~l178;
assign a8092 = a8090 & ~l176;
assign a8094 = a8092 & l174;
assign a8096 = ~a8094 & a8086;
assign a8098 = a8096 & a8082;
assign a8100 = a8082 & l210;
assign a8102 = a8100 & a7932;
assign a8104 = a8102 & ~a8094;
assign a8106 = a8104 & l172;
assign a8108 = a8106 & l170;
assign a8110 = a8108 & ~l168;
assign a8112 = a8110 & ~l166;
assign a8114 = a8112 & l164;
assign a8116 = a8084 & a7960;
assign a8118 = a8116 & ~a8094;
assign a8120 = a8118 & l172;
assign a8122 = a8120 & l170;
assign a8124 = a8122 & ~l168;
assign a8126 = a8124 & ~l166;
assign a8128 = a8126 & l164;
assign a8130 = a8100 & a7960;
assign a8132 = a8130 & ~a8094;
assign a8134 = a8132 & l172;
assign a8136 = a8134 & l170;
assign a8138 = a8136 & ~l168;
assign a8140 = a8138 & ~l166;
assign a8142 = a8140 & l164;
assign a8144 = a8082 & a7938;
assign a8146 = a8144 & l194;
assign a8148 = a8146 & ~a8094;
assign a8150 = a8148 & l172;
assign a8152 = a8150 & l170;
assign a8154 = a8152 & ~l168;
assign a8156 = a8154 & ~l166;
assign a8158 = a8156 & l164;
assign a8160 = a8082 & ~a7950;
assign a8162 = a8160 & l204;
assign a8164 = a8162 & ~a8094;
assign a8166 = a8164 & l172;
assign a8168 = a8166 & l170;
assign a8170 = a8168 & ~l168;
assign a8172 = a8170 & ~l166;
assign a8174 = a8172 & l164;
assign a8176 = a8082 & ~l208;
assign a8178 = a8176 & l224;
assign a8180 = a8178 & l198;
assign a8182 = a8180 & ~a8094;
assign a8184 = a8182 & l172;
assign a8186 = a8184 & l170;
assign a8188 = a8186 & ~l168;
assign a8190 = a8188 & ~l166;
assign a8192 = a8190 & l164;
assign a8194 = a8082 & l208;
assign a8196 = a8194 & a7950;
assign a8198 = a8196 & l186;
assign a8200 = a8198 & ~l194;
assign a8202 = a8200 & ~a8094;
assign a8204 = a8202 & a8082;
assign a8206 = a8194 & l210;
assign a8208 = a8206 & l214;
assign a8210 = a8208 & a7960;
assign a8212 = a8210 & l186;
assign a8214 = a8212 & ~l194;
assign a8216 = a8214 & ~a8094;
assign a8218 = a8216 & l172;
assign a8220 = a8218 & l170;
assign a8222 = a8220 & ~l168;
assign a8224 = a8222 & ~l166;
assign a8226 = a8224 & l164;
assign a8228 = a8082 & ~l210;
assign a8230 = a8228 & a7924;
assign a8232 = a8230 & l186;
assign a8234 = a8232 & ~l194;
assign a8236 = a8234 & ~a8094;
assign a8238 = a8236 & l172;
assign a8240 = a8238 & l170;
assign a8242 = a8240 & ~l168;
assign a8244 = a8242 & ~l166;
assign a8246 = a8244 & l164;
assign a8248 = a8100 & a7924;
assign a8250 = a8248 & l186;
assign a8252 = a8250 & ~l194;
assign a8254 = a8252 & ~a8094;
assign a8256 = a8254 & l172;
assign a8258 = a8256 & l170;
assign a8260 = a8258 & ~l168;
assign a8262 = a8260 & ~l166;
assign a8264 = a8262 & l164;
assign a8266 = a8100 & l214;
assign a8268 = a8266 & a7932;
assign a8270 = a8268 & l186;
assign a8272 = a8270 & ~l194;
assign a8274 = a8272 & ~a8094;
assign a8276 = a8274 & l172;
assign a8278 = a8276 & l170;
assign a8280 = a8278 & ~l168;
assign a8282 = a8280 & ~l166;
assign a8284 = a8282 & l164;
assign a8286 = a8144 & l186;
assign a8288 = a8286 & ~l194;
assign a8290 = a8288 & ~a8094;
assign a8292 = a8290 & l172;
assign a8294 = a8292 & l170;
assign a8296 = a8294 & ~l168;
assign a8298 = a8296 & ~l166;
assign a8300 = a8298 & l164;
assign a8302 = a8176 & a7950;
assign a8304 = a8302 & l186;
assign a8306 = a8304 & ~l194;
assign a8308 = a8306 & ~a8094;
assign a8310 = a8308 & l172;
assign a8312 = a8310 & l170;
assign a8314 = a8312 & ~l168;
assign a8316 = a8314 & ~l166;
assign a8318 = a8316 & l164;
assign a8320 = a8176 & l210;
assign a8322 = a8320 & l214;
assign a8324 = a8322 & a7960;
assign a8326 = a8324 & l186;
assign a8328 = a8326 & ~l194;
assign a8330 = a8328 & ~a8094;
assign a8332 = a8330 & l172;
assign a8334 = a8332 & l170;
assign a8336 = a8334 & ~l168;
assign a8338 = a8336 & ~l166;
assign a8340 = a8338 & l164;
assign a8342 = a8082 & l200;
assign a8344 = a8342 & ~a8094;
assign a8346 = a8344 & l172;
assign a8348 = a8346 & l170;
assign a8350 = a8348 & ~l168;
assign a8352 = a8350 & ~l166;
assign a8354 = a8352 & l164;
assign a8356 = a8082 & ~l186;
assign a8358 = a8356 & ~a8094;
assign a8360 = a8358 & l172;
assign a8362 = a8360 & l170;
assign a8364 = a8362 & ~l168;
assign a8366 = a8364 & ~l166;
assign a8368 = a8366 & l164;
assign a8370 = a8082 & a7950;
assign a8372 = a8370 & l222;
assign a8374 = a8372 & l186;
assign a8376 = a8374 & l198;
assign a8378 = a8376 & ~a8094;
assign a8380 = a8378 & l172;
assign a8382 = a8380 & l170;
assign a8384 = a8382 & ~l168;
assign a8386 = a8384 & ~l166;
assign a8388 = a8386 & l164;
assign a8390 = a8198 & l198;
assign a8392 = a8390 & ~a8094;
assign a8394 = a8392 & l172;
assign a8396 = a8394 & l170;
assign a8398 = a8396 & ~l168;
assign a8400 = a8398 & ~l166;
assign a8402 = a8400 & l164;
assign a8404 = a8266 & a7960;
assign a8406 = a8404 & l222;
assign a8408 = a8406 & l186;
assign a8410 = a8408 & l198;
assign a8412 = a8410 & ~a8094;
assign a8414 = a8412 & l172;
assign a8416 = a8414 & l170;
assign a8418 = a8416 & ~l168;
assign a8420 = a8418 & ~l166;
assign a8422 = a8420 & l164;
assign a8424 = a8212 & l198;
assign a8426 = a8424 & ~a8094;
assign a8428 = a8426 & l172;
assign a8430 = a8428 & l170;
assign a8432 = a8430 & ~l168;
assign a8434 = a8432 & ~l166;
assign a8436 = a8434 & l164;
assign a8438 = a8230 & l222;
assign a8440 = a8438 & l186;
assign a8442 = a8440 & l198;
assign a8444 = a8442 & ~a8094;
assign a8446 = a8444 & l172;
assign a8448 = a8446 & l170;
assign a8450 = a8448 & ~l168;
assign a8452 = a8450 & ~l166;
assign a8454 = a8452 & l164;
assign a8456 = a8194 & ~l210;
assign a8458 = a8456 & a7924;
assign a8460 = a8458 & l186;
assign a8462 = a8460 & l198;
assign a8464 = a8462 & ~a8094;
assign a8466 = a8464 & l172;
assign a8468 = a8466 & l170;
assign a8470 = a8468 & ~l168;
assign a8472 = a8470 & ~l166;
assign a8474 = a8472 & l164;
assign a8476 = a8248 & l222;
assign a8478 = a8476 & l186;
assign a8480 = a8478 & l198;
assign a8482 = a8480 & ~a8094;
assign a8484 = a8482 & l172;
assign a8486 = a8484 & l170;
assign a8488 = a8486 & ~l168;
assign a8490 = a8488 & ~l166;
assign a8492 = a8490 & l164;
assign a8494 = a8206 & a7924;
assign a8496 = a8494 & l186;
assign a8498 = a8496 & l198;
assign a8500 = a8498 & ~a8094;
assign a8502 = a8500 & l172;
assign a8504 = a8502 & l170;
assign a8506 = a8504 & ~l168;
assign a8508 = a8506 & ~l166;
assign a8510 = a8508 & l164;
assign a8512 = a8268 & l222;
assign a8514 = a8512 & l186;
assign a8516 = a8514 & l198;
assign a8518 = a8516 & ~a8094;
assign a8520 = a8518 & l172;
assign a8522 = a8520 & l170;
assign a8524 = a8522 & ~l168;
assign a8526 = a8524 & ~l166;
assign a8528 = a8526 & l164;
assign a8530 = a8208 & a7932;
assign a8532 = a8530 & l186;
assign a8534 = a8532 & l198;
assign a8536 = a8534 & ~a8094;
assign a8538 = a8536 & l172;
assign a8540 = a8538 & l170;
assign a8542 = a8540 & ~l168;
assign a8544 = a8542 & ~l166;
assign a8546 = a8544 & l164;
assign a8548 = a6722 & l166;
assign a8550 = a8548 & ~l164;
assign a8552 = a8550 & l216;
assign a8554 = a8552 & ~l226;
assign a8556 = a8554 & i54;
assign a8558 = a8550 & l236;
assign a8560 = a8558 & ~i64;
assign a8562 = a8548 & l234;
assign a8564 = a8562 & ~i62;
assign a8566 = a8550 & ~a7924;
assign a8568 = a8566 & ~i74;
assign a8570 = a8568 & ~i72;
assign a8572 = a8570 & ~i70;
assign a8574 = a8550 & ~a7932;
assign a8576 = a8574 & i74;
assign a8578 = a8576 & ~i72;
assign a8580 = a8578 & ~i70;
assign a8582 = a8550 & ~a7938;
assign a8584 = a8582 & ~i70;
assign a8586 = a8584 & ~i74;
assign a8588 = a8586 & i72;
assign a8590 = a8550 & ~a7960;
assign a8592 = a8590 & ~i74;
assign a8594 = a8592 & ~i72;
assign a8596 = a8594 & i70;
assign a8598 = a8550 & l186;
assign a8600 = a8598 & ~i14;
assign a8602 = a8550 & ~l198;
assign a8604 = a8602 & i26;
assign a8606 = a8550 & ~l200;
assign a8608 = a8606 & i28;
assign a8610 = a8550 & ~l204;
assign a8612 = a8610 & i32;
assign a8614 = a8550 & ~l206;
assign a8616 = a8614 & i34;
assign a8618 = a8548 & ~l216;
assign a8620 = a8618 & l208;
assign a8622 = a8620 & ~i36;
assign a8624 = a7860 & l166;
assign a8626 = a8624 & ~l164;
assign a8628 = a8626 & l236;
assign a8630 = a8628 & ~i64;
assign a8632 = a8626 & l216;
assign a8634 = a8632 & ~l226;
assign a8636 = a8634 & i54;
assign a8638 = a8626 & ~l210;
assign a8640 = a8638 & i38;
assign a8642 = a8640 & l214;
assign a8644 = a8642 & ~l228;
assign a8646 = a8626 & l214;
assign a8648 = a8646 & ~i42;
assign a8650 = a8626 & ~l204;
assign a8652 = a8650 & i32;
assign a8654 = a8624 & l234;
assign a8656 = a8654 & ~i62;
assign a8658 = a8626 & ~a7924;
assign a8660 = a8658 & ~i74;
assign a8662 = a8660 & ~i72;
assign a8664 = a8662 & ~i70;
assign a8666 = a8626 & ~a7932;
assign a8668 = a8666 & i74;
assign a8670 = a8668 & ~i72;
assign a8672 = a8670 & ~i70;
assign a8674 = a8626 & ~a7938;
assign a8676 = a8674 & ~i70;
assign a8678 = a8676 & ~i74;
assign a8680 = a8678 & i72;
assign a8682 = a8626 & ~a7950;
assign a8684 = a8682 & i74;
assign a8686 = a8684 & i72;
assign a8688 = a8686 & ~i70;
assign a8690 = a8626 & l186;
assign a8692 = a8690 & ~i14;
assign a8694 = a8626 & ~l200;
assign a8696 = a8694 & i28;
assign a8698 = a8626 & ~l198;
assign a8700 = a8698 & i26;
assign a8702 = a8624 & ~l216;
assign a8704 = a8702 & l208;
assign a8706 = a8704 & ~i36;
assign a8708 = a6726 & l236;
assign a8710 = a8708 & ~i64;
assign a8712 = a6726 & l216;
assign a8714 = a8712 & ~l226;
assign a8716 = a8714 & i54;
assign a8718 = a6726 & ~l204;
assign a8720 = a8718 & i32;
assign a8722 = a6724 & l234;
assign a8724 = a8722 & ~i62;
assign a8726 = ~a7932 & a6726;
assign a8728 = a8726 & i74;
assign a8730 = a8728 & ~i72;
assign a8732 = a8730 & ~i70;
assign a8734 = ~a7938 & a6726;
assign a8736 = a8734 & ~i70;
assign a8738 = a8736 & ~i74;
assign a8740 = a8738 & i72;
assign a8742 = ~a7950 & a6726;
assign a8744 = a8742 & i74;
assign a8746 = a8744 & i72;
assign a8748 = a8746 & ~i70;
assign a8750 = ~a7960 & a6726;
assign a8752 = a8750 & ~i74;
assign a8754 = a8752 & ~i72;
assign a8756 = a8754 & i70;
assign a8758 = a6726 & l186;
assign a8760 = a8758 & ~i14;
assign a8762 = a6726 & ~l200;
assign a8764 = a8762 & i28;
assign a8766 = a6726 & ~l198;
assign a8768 = a8766 & i26;
assign a8770 = a6724 & ~l210;
assign a8772 = a8770 & i38;
assign a8774 = a8772 & ~l228;
assign a8776 = a7862 & ~l164;
assign a8778 = a8776 & l236;
assign a8780 = a8778 & ~i64;
assign a8782 = a8776 & l216;
assign a8784 = a8782 & ~l226;
assign a8786 = a8784 & i54;
assign a8788 = a8776 & ~l204;
assign a8790 = a8788 & i32;
assign a8792 = a7862 & l234;
assign a8794 = a8792 & ~i62;
assign a8796 = a8776 & ~a7932;
assign a8798 = a8796 & i74;
assign a8800 = a8798 & ~i72;
assign a8802 = a8800 & ~i70;
assign a8804 = a8776 & ~a7938;
assign a8806 = a8804 & ~i70;
assign a8808 = a8806 & ~i74;
assign a8810 = a8808 & i72;
assign a8812 = a8776 & ~a7950;
assign a8814 = a8812 & i74;
assign a8816 = a8814 & i72;
assign a8818 = a8816 & ~i70;
assign a8820 = a8776 & ~a7960;
assign a8822 = a8820 & ~i74;
assign a8824 = a8822 & ~i72;
assign a8826 = a8824 & i70;
assign a8828 = a8776 & l186;
assign a8830 = a8828 & ~i14;
assign a8832 = a8776 & ~l198;
assign a8834 = a8832 & i26;
assign a8836 = a8776 & ~l200;
assign a8838 = a8836 & i28;
assign a8840 = a7862 & ~l220;
assign a8842 = a8840 & i48;
assign a8844 = a8006 & ~l166;
assign a8846 = a8844 & ~l164;
assign a8848 = a8846 & l236;
assign a8850 = a8848 & ~i64;
assign a8852 = a8846 & l216;
assign a8854 = a8852 & ~l226;
assign a8856 = a8854 & i54;
assign a8858 = a8846 & l214;
assign a8860 = a8858 & ~i42;
assign a8862 = a8846 & ~l210;
assign a8864 = a8862 & i38;
assign a8866 = a8864 & l214;
assign a8868 = a8866 & ~l228;
assign a8870 = a8846 & ~l204;
assign a8872 = a8870 & i32;
assign a8874 = a8844 & l234;
assign a8876 = a8874 & ~i62;
assign a8878 = a8846 & ~a7924;
assign a8880 = a8878 & ~i74;
assign a8882 = a8880 & ~i72;
assign a8884 = a8882 & ~i70;
assign a8886 = a8846 & ~a7938;
assign a8888 = a8886 & ~i70;
assign a8890 = a8888 & ~i74;
assign a8892 = a8890 & i72;
assign a8894 = a8846 & ~a7950;
assign a8896 = a8894 & i74;
assign a8898 = a8896 & i72;
assign a8900 = a8898 & ~i70;
assign a8902 = a8846 & ~a7960;
assign a8904 = a8902 & ~i74;
assign a8906 = a8904 & ~i72;
assign a8908 = a8906 & i70;
assign a8910 = a8846 & l186;
assign a8912 = a8910 & ~i14;
assign a8914 = a8846 & ~l200;
assign a8916 = a8914 & i28;
assign a8918 = a8846 & ~l198;
assign a8920 = a8918 & i26;
assign a8922 = a8844 & ~l220;
assign a8924 = a8922 & i48;
assign a8926 = ~l172 & l170;
assign a8928 = a8926 & l168;
assign a8930 = a8928 & ~l166;
assign a8932 = a8930 & ~l164;
assign a8934 = a8932 & l236;
assign a8936 = a8934 & ~i64;
assign a8938 = a8932 & ~l204;
assign a8940 = a8938 & i32;
assign a8942 = a8932 & ~l206;
assign a8944 = a8942 & i34;
assign a8946 = a8932 & ~l198;
assign a8948 = a8946 & i26;
assign a8950 = a8930 & l234;
assign a8952 = a8950 & ~i62;
assign a8954 = a8932 & ~a7924;
assign a8956 = a8954 & ~i74;
assign a8958 = a8956 & ~i72;
assign a8960 = a8958 & ~i70;
assign a8962 = a8932 & ~a7932;
assign a8964 = a8962 & i74;
assign a8966 = a8964 & ~i72;
assign a8968 = a8966 & ~i70;
assign a8970 = a8932 & ~a7950;
assign a8972 = a8970 & i74;
assign a8974 = a8972 & i72;
assign a8976 = a8974 & ~i70;
assign a8978 = a8932 & ~a7960;
assign a8980 = a8978 & ~i74;
assign a8982 = a8980 & ~i72;
assign a8984 = a8982 & i70;
assign a8986 = a8932 & l186;
assign a8988 = a8986 & ~i14;
assign a8990 = a8932 & ~l200;
assign a8992 = a8990 & i28;
assign a8994 = a6720 & l168;
assign a8996 = a8994 & ~l166;
assign a8998 = a8996 & ~l164;
assign a9000 = a8998 & l236;
assign a9002 = a9000 & ~i64;
assign a9004 = a8998 & l216;
assign a9006 = a9004 & ~l226;
assign a9008 = a9006 & i54;
assign a9010 = a8996 & l234;
assign a9012 = a9010 & ~i62;
assign a9014 = a8998 & ~a7924;
assign a9016 = a9014 & ~i74;
assign a9018 = a9016 & ~i72;
assign a9020 = a9018 & ~i70;
assign a9022 = a8998 & ~a7932;
assign a9024 = a9022 & i74;
assign a9026 = a9024 & ~i72;
assign a9028 = a9026 & ~i70;
assign a9030 = a8998 & ~a7938;
assign a9032 = a9030 & ~i70;
assign a9034 = a9032 & ~i74;
assign a9036 = a9034 & i72;
assign a9038 = a8998 & ~a7960;
assign a9040 = a9038 & ~i74;
assign a9042 = a9040 & ~i72;
assign a9044 = a9042 & i70;
assign a9046 = a8998 & l186;
assign a9048 = a9046 & ~i14;
assign a9050 = a8998 & ~l198;
assign a9052 = a9050 & i26;
assign a9054 = a8998 & ~l200;
assign a9056 = a9054 & i28;
assign a9058 = a8998 & ~l204;
assign a9060 = a9058 & i32;
assign a9062 = a8996 & ~l220;
assign a9064 = a9062 & i48;
assign a9066 = a7858 & ~l168;
assign a9068 = a9066 & l166;
assign a9070 = a9068 & ~l164;
assign a9072 = a9070 & l236;
assign a9074 = a9072 & ~i64;
assign a9076 = a9070 & l216;
assign a9078 = a9076 & ~l226;
assign a9080 = a9078 & i54;
assign a9082 = a9070 & l214;
assign a9084 = a9082 & ~i42;
assign a9086 = a9070 & ~l210;
assign a9088 = a9086 & i38;
assign a9090 = a9088 & l214;
assign a9092 = a9090 & ~l228;
assign a9094 = a9070 & ~l204;
assign a9096 = a9094 & i32;
assign a9098 = a9068 & l234;
assign a9100 = a9098 & ~i62;
assign a9102 = a9070 & ~a7924;
assign a9104 = a9102 & ~i74;
assign a9106 = a9104 & ~i72;
assign a9108 = a9106 & ~i70;
assign a9110 = a9070 & ~a7932;
assign a9112 = a9110 & i74;
assign a9114 = a9112 & ~i72;
assign a9116 = a9114 & ~i70;
assign a9118 = a9070 & ~a7938;
assign a9120 = a9118 & ~i70;
assign a9122 = a9120 & ~i74;
assign a9124 = a9122 & i72;
assign a9126 = a9070 & ~a7950;
assign a9128 = a9126 & i74;
assign a9130 = a9128 & i72;
assign a9132 = a9130 & ~i70;
assign a9134 = a9070 & l186;
assign a9136 = a9134 & ~i14;
assign a9138 = a9070 & ~l200;
assign a9140 = a9138 & i28;
assign a9142 = a9070 & ~l198;
assign a9144 = a9142 & i26;
assign a9146 = a9068 & ~l220;
assign a9148 = a9146 & i48;
assign a9150 = a8926 & ~l168;
assign a9152 = a9150 & ~l166;
assign a9154 = a9152 & ~l164;
assign a9156 = a9154 & l236;
assign a9158 = a9156 & ~i64;
assign a9160 = a9152 & l234;
assign a9162 = a9160 & ~i62;
assign a9164 = a9154 & ~l198;
assign a9166 = a9164 & i26;
assign a9168 = a9154 & ~l202;
assign a9170 = a9168 & i30;
assign a9172 = a9154 & ~l204;
assign a9174 = a9172 & i32;
assign a9176 = a9154 & ~l206;
assign a9178 = a9176 & i34;
assign a9180 = a9154 & ~l196;
assign a9182 = a9180 & i24;
assign a9184 = a9066 & ~l166;
assign a9186 = a9184 & ~l164;
assign a9188 = a9186 & l236;
assign a9190 = a9188 & ~i64;
assign a9192 = a9186 & ~l240;
assign a9194 = a9192 & i68;
assign a9196 = a9184 & ~l196;
assign a9198 = a9196 & i24;
assign a9200 = a9186 & ~a7924;
assign a9202 = a9200 & ~i74;
assign a9204 = a9202 & ~i72;
assign a9206 = a9204 & ~i70;
assign a9208 = a9186 & ~a7932;
assign a9210 = a9208 & i74;
assign a9212 = a9210 & ~i72;
assign a9214 = a9212 & ~i70;
assign a9216 = a9186 & ~a7938;
assign a9218 = a9216 & ~i70;
assign a9220 = a9218 & ~i74;
assign a9222 = a9220 & i72;
assign a9224 = a9186 & ~a7950;
assign a9226 = a9224 & i74;
assign a9228 = a9226 & i72;
assign a9230 = a9228 & ~i70;
assign a9232 = a9186 & ~a7960;
assign a9234 = a9232 & ~i74;
assign a9236 = a9234 & ~i72;
assign a9238 = a9236 & i70;
assign a9240 = a8004 & ~l168;
assign a9242 = a9240 & l166;
assign a9244 = a9242 & ~l164;
assign a9246 = a9244 & l236;
assign a9248 = a9246 & ~i64;
assign a9250 = a9244 & l186;
assign a9252 = a9250 & ~i14;
assign a9254 = a9244 & ~l198;
assign a9256 = a9254 & i26;
assign a9258 = a9242 & l240;
assign a9260 = a9258 & ~i68;
assign a9262 = a9244 & ~a7924;
assign a9264 = a9262 & ~i74;
assign a9266 = a9264 & ~i72;
assign a9268 = a9266 & ~i70;
assign a9270 = a9244 & ~a7932;
assign a9272 = a9270 & i74;
assign a9274 = a9272 & ~i72;
assign a9276 = a9274 & ~i70;
assign a9278 = a9244 & ~a7938;
assign a9280 = a9278 & ~i70;
assign a9282 = a9280 & ~i74;
assign a9284 = a9282 & i72;
assign a9286 = a9244 & ~a7950;
assign a9288 = a9286 & i74;
assign a9290 = a9288 & i72;
assign a9292 = a9290 & ~i70;
assign a9294 = a9244 & ~a7960;
assign a9296 = a9294 & ~i74;
assign a9298 = a9296 & ~i72;
assign a9300 = a9298 & i70;
assign a9302 = a9240 & ~l166;
assign a9304 = a9302 & ~l164;
assign a9306 = a9304 & l236;
assign a9308 = a9306 & ~i64;
assign a9310 = a9302 & ~l240;
assign a9312 = a9310 & i68;
assign a9314 = a9304 & ~a7924;
assign a9316 = a9314 & ~i74;
assign a9318 = a9316 & ~i72;
assign a9320 = a9318 & ~i70;
assign a9322 = a9304 & ~a7932;
assign a9324 = a9322 & i74;
assign a9326 = a9324 & ~i72;
assign a9328 = a9326 & ~i70;
assign a9330 = a9304 & ~a7938;
assign a9332 = a9330 & ~i70;
assign a9334 = a9332 & ~i74;
assign a9336 = a9334 & i72;
assign a9338 = a9304 & ~a7950;
assign a9340 = a9338 & i74;
assign a9342 = a9340 & i72;
assign a9344 = a9342 & ~i70;
assign a9346 = a9304 & ~a7960;
assign a9348 = a9346 & ~i74;
assign a9350 = a9348 & ~i72;
assign a9352 = a9350 & i70;
assign a9354 = a9302 & l164;
assign a9356 = a9354 & l236;
assign a9358 = a9356 & ~i64;
assign a9360 = a9354 & l216;
assign a9362 = a9360 & ~l226;
assign a9364 = a9362 & i54;
assign a9366 = a9354 & l186;
assign a9368 = a9366 & ~i14;
assign a9370 = a9354 & l208;
assign a9372 = a9370 & ~i36;
assign a9374 = a9354 & l234;
assign a9376 = a9374 & ~i62;
assign a9378 = a9354 & ~a7924;
assign a9380 = a9378 & ~i74;
assign a9382 = a9380 & ~i72;
assign a9384 = a9382 & ~i70;
assign a9386 = a9354 & ~a7932;
assign a9388 = a9386 & i74;
assign a9390 = a9388 & ~i72;
assign a9392 = a9390 & ~i70;
assign a9394 = a9354 & ~a7938;
assign a9396 = a9394 & ~i70;
assign a9398 = a9396 & ~i74;
assign a9400 = a9398 & i72;
assign a9402 = a9354 & ~a7960;
assign a9404 = a9402 & ~i74;
assign a9406 = a9404 & ~i72;
assign a9408 = a9406 & i70;
assign a9410 = a9354 & ~l200;
assign a9412 = a9410 & i28;
assign a9414 = a9354 & ~l202;
assign a9416 = a9414 & i30;
assign a9418 = a9354 & ~l204;
assign a9420 = a9418 & i32;
assign a9422 = a9354 & ~l206;
assign a9424 = a9422 & i34;
assign a9426 = a9354 & ~l196;
assign a9428 = a9426 & i24;
assign a9430 = a9354 & ~l212;
assign a9432 = a9430 & i40;
assign a9434 = a9354 & l210;
assign a9436 = a9434 & ~i38;
assign a9438 = a9354 & ~l210;
assign a9440 = a9438 & i38;
assign a9442 = a9440 & ~l228;
assign a9444 = a9354 & ~l214;
assign a9446 = a9444 & i42;
assign a9448 = a9446 & ~l228;
assign a9450 = a9354 & l214;
assign a9452 = a9450 & ~i42;
assign a9454 = a9354 & ~l220;
assign a9456 = a9454 & i48;
assign a9458 = a9152 & l164;
assign a9460 = a9458 & l236;
assign a9462 = a9460 & ~i64;
assign a9464 = a9458 & l216;
assign a9466 = a9464 & ~l226;
assign a9468 = a9466 & i54;
assign a9470 = a9458 & l214;
assign a9472 = a9470 & ~i42;
assign a9474 = a9458 & ~l210;
assign a9476 = a9474 & i38;
assign a9478 = a9476 & l214;
assign a9480 = a9478 & ~l228;
assign a9482 = a9458 & l208;
assign a9484 = a9482 & ~i36;
assign a9486 = a9458 & l186;
assign a9488 = a9486 & ~i14;
assign a9490 = a9458 & l234;
assign a9492 = a9490 & ~i62;
assign a9494 = a9458 & ~a7924;
assign a9496 = a9494 & ~i74;
assign a9498 = a9496 & ~i72;
assign a9500 = a9498 & ~i70;
assign a9502 = a9458 & ~a7932;
assign a9504 = a9502 & i74;
assign a9506 = a9504 & ~i72;
assign a9508 = a9506 & ~i70;
assign a9510 = a9458 & ~a7938;
assign a9512 = a9510 & ~i70;
assign a9514 = a9512 & ~i74;
assign a9516 = a9514 & i72;
assign a9518 = a9458 & ~a7950;
assign a9520 = a9518 & i74;
assign a9522 = a9520 & i72;
assign a9524 = a9522 & ~i70;
assign a9526 = a9458 & ~l200;
assign a9528 = a9526 & i28;
assign a9530 = a9458 & ~l202;
assign a9532 = a9530 & i30;
assign a9534 = a9458 & ~l204;
assign a9536 = a9534 & i32;
assign a9538 = a9458 & ~l206;
assign a9540 = a9538 & i34;
assign a9542 = a9458 & ~l196;
assign a9544 = a9542 & i24;
assign a9546 = a9458 & ~l212;
assign a9548 = a9546 & i40;
assign a9550 = a9458 & ~l220;
assign a9552 = a9550 & i48;
assign a9554 = a8928 & l166;
assign a9556 = a9554 & ~l164;
assign a9558 = a9556 & l236;
assign a9560 = a9558 & ~i64;
assign a9562 = a9556 & l216;
assign a9564 = a9562 & ~l226;
assign a9566 = a9564 & i54;
assign a9568 = a9556 & l186;
assign a9570 = a9568 & ~i14;
assign a9572 = a9556 & l234;
assign a9574 = a9572 & ~i62;
assign a9576 = a9556 & ~a7932;
assign a9578 = a9576 & i74;
assign a9580 = a9578 & ~i72;
assign a9582 = a9580 & ~i70;
assign a9584 = a9556 & ~a7938;
assign a9586 = a9584 & ~i70;
assign a9588 = a9586 & ~i74;
assign a9590 = a9588 & i72;
assign a9592 = a9556 & ~a7950;
assign a9594 = a9592 & i74;
assign a9596 = a9594 & i72;
assign a9598 = a9596 & ~i70;
assign a9600 = a9556 & ~a7960;
assign a9602 = a9600 & ~i74;
assign a9604 = a9602 & ~i72;
assign a9606 = a9604 & i70;
assign a9608 = a9556 & ~l200;
assign a9610 = a9608 & i28;
assign a9612 = a9556 & ~l202;
assign a9614 = a9612 & i30;
assign a9616 = a9556 & ~l204;
assign a9618 = a9616 & i32;
assign a9620 = a9556 & ~l206;
assign a9622 = a9620 & i34;
assign a9624 = a9556 & ~l196;
assign a9626 = a9624 & i24;
assign a9628 = a9554 & ~l210;
assign a9630 = a9628 & i38;
assign a9632 = a9630 & ~l228;
assign a9634 = a8994 & l166;
assign a9636 = a9634 & ~l164;
assign a9638 = a9636 & l236;
assign a9640 = a9638 & ~i64;
assign a9642 = a9636 & l216;
assign a9644 = a9642 & ~l226;
assign a9646 = a9644 & i54;
assign a9648 = a9636 & l186;
assign a9650 = a9648 & ~i14;
assign a9652 = a9636 & l234;
assign a9654 = a9652 & ~i62;
assign a9656 = a9636 & ~a7932;
assign a9658 = a9656 & i74;
assign a9660 = a9658 & ~i72;
assign a9662 = a9660 & ~i70;
assign a9664 = a9636 & ~a7938;
assign a9666 = a9664 & ~i70;
assign a9668 = a9666 & ~i74;
assign a9670 = a9668 & i72;
assign a9672 = a9636 & ~a7950;
assign a9674 = a9672 & i74;
assign a9676 = a9674 & i72;
assign a9678 = a9676 & ~i70;
assign a9680 = a9636 & ~a7960;
assign a9682 = a9680 & ~i74;
assign a9684 = a9682 & ~i72;
assign a9686 = a9684 & i70;
assign a9688 = a9636 & ~l200;
assign a9690 = a9688 & i28;
assign a9692 = a9636 & ~l202;
assign a9694 = a9692 & i30;
assign a9696 = a9636 & ~l204;
assign a9698 = a9696 & i32;
assign a9700 = a9636 & ~l206;
assign a9702 = a9700 & i34;
assign a9704 = a9636 & ~l196;
assign a9706 = a9704 & i24;
assign a9708 = a9634 & l214;
assign a9710 = a9708 & ~i42;
assign a9712 = ~l172 & ~l168;
assign a9714 = ~l170 & ~l166;
assign a9716 = a9714 & l164;
assign a9718 = a9716 & ~l220;
assign a9720 = a9718 & i48;
assign a9722 = l236 & ~i64;
assign a9724 = a9150 & l166;
assign a9726 = a9724 & l234;
assign a9728 = a9726 & ~i62;
assign a9730 = ~l206 & i34;
assign a9732 = ~l196 & i24;
assign a9734 = ~l202 & i30;
assign a9736 = ~l200 & i28;
assign a9738 = ~l198 & i26;
assign a9740 = l186 & ~i14;
assign a9742 = ~a7960 & a358;
assign a9744 = a7944 & ~a7938;
assign a9746 = ~a7932 & a354;
assign a9748 = a7928 & ~a7924;
assign a9750 = ~a9748 & ~a9746;
assign a9752 = a9750 & ~a9744;
assign a9754 = a9752 & ~a9742;
assign a9756 = a9754 & ~a9740;
assign a9758 = a9756 & ~a9738;
assign a9760 = a9758 & ~a9736;
assign a9762 = a9760 & ~a9734;
assign a9764 = a9762 & ~a9732;
assign a9766 = a9764 & ~a9730;
assign a9768 = ~a9766 & ~a9728;
assign a9770 = ~a9768 & ~a9722;
assign a9772 = l170 & l166;
assign a9774 = a9772 & ~l164;
assign a9776 = a9774 & ~a9770;
assign a9778 = a9716 & ~l212;
assign a9780 = a9778 & i40;
assign a9782 = a9716 & ~l196;
assign a9784 = a9782 & i24;
assign a9786 = a9716 & ~l206;
assign a9788 = a9786 & i34;
assign a9790 = a9716 & ~l204;
assign a9792 = a9790 & i32;
assign a9794 = a9716 & ~l202;
assign a9796 = a9794 & i30;
assign a9798 = a9716 & ~l200;
assign a9800 = a9798 & i28;
assign a9802 = a9716 & ~a7960;
assign a9804 = a9802 & ~i74;
assign a9806 = a9804 & ~i72;
assign a9808 = a9806 & i70;
assign a9810 = a9716 & ~a7950;
assign a9812 = a9810 & i74;
assign a9814 = a9812 & i72;
assign a9816 = a9814 & ~i70;
assign a9818 = a9716 & ~a7938;
assign a9820 = a9818 & ~i70;
assign a9822 = a9820 & ~i74;
assign a9824 = a9822 & i72;
assign a9826 = a9716 & ~a7924;
assign a9828 = a9826 & ~i74;
assign a9830 = a9828 & ~i72;
assign a9832 = a9830 & ~i70;
assign a9834 = a9716 & l234;
assign a9836 = a9834 & ~i62;
assign a9838 = a9716 & l186;
assign a9840 = a9838 & ~i14;
assign a9842 = a9716 & ~l210;
assign a9844 = a9842 & i38;
assign a9846 = a9844 & l214;
assign a9848 = a9846 & ~l228;
assign a9850 = a9716 & l214;
assign a9852 = a9850 & ~i42;
assign a9854 = a9716 & l216;
assign a9856 = a9854 & ~l226;
assign a9858 = a9856 & i54;
assign a9860 = a9716 & l236;
assign a9862 = a9860 & ~i64;
assign a9864 = ~a9862 & ~a9858;
assign a9866 = a9864 & ~a9852;
assign a9868 = a9866 & ~a9848;
assign a9870 = a9868 & ~a9840;
assign a9872 = a9870 & ~a9836;
assign a9874 = a9872 & ~a9832;
assign a9876 = a9874 & ~a9824;
assign a9878 = a9876 & ~a9816;
assign a9880 = a9878 & ~a9808;
assign a9882 = a9880 & ~a9800;
assign a9884 = a9882 & ~a9796;
assign a9886 = a9884 & ~a9792;
assign a9888 = a9886 & ~a9788;
assign a9890 = a9888 & ~a9784;
assign a9892 = a9890 & ~a9780;
assign a9894 = a9892 & ~a9776;
assign a9896 = a9894 & ~a9720;
assign a9898 = a9634 & l210;
assign a9900 = a9898 & ~l214;
assign a9902 = a9900 & i42;
assign a9904 = a9902 & ~l228;
assign a9906 = a9634 & ~l220;
assign a9908 = a9906 & i48;
assign a9910 = a9898 & ~i38;
assign a9912 = ~a9910 & ~a9908;
assign a9914 = a9912 & ~a9904;
assign a9916 = a9914 & ~a9896;
assign a9918 = a9916 & a9712;
assign a9920 = a9918 & ~a9710;
assign a9922 = ~a9920 & ~a9706;
assign a9924 = a9922 & ~a9702;
assign a9926 = a9924 & ~a9698;
assign a9928 = a9926 & ~a9694;
assign a9930 = a9928 & ~a9690;
assign a9932 = a9930 & ~a9686;
assign a9934 = a9932 & ~a9678;
assign a9936 = a9934 & ~a9670;
assign a9938 = a9936 & ~a9662;
assign a9940 = a9938 & ~a9654;
assign a9942 = a9940 & ~a9650;
assign a9944 = a9942 & ~a9646;
assign a9946 = a9944 & ~a9640;
assign a9948 = a9554 & ~l220;
assign a9950 = a9948 & i48;
assign a9952 = a9554 & ~l218;
assign a9954 = a9952 & i46;
assign a9956 = a9554 & ~l212;
assign a9958 = a9956 & i40;
assign a9960 = a9554 & l214;
assign a9962 = a9960 & ~i42;
assign a9964 = a9628 & ~l214;
assign a9966 = a9964 & i42;
assign a9968 = a9966 & ~l228;
assign a9970 = ~a9968 & ~a9962;
assign a9972 = a9970 & ~a9958;
assign a9974 = a9972 & ~a9954;
assign a9976 = a9974 & ~a9950;
assign a9978 = a9976 & ~a9946;
assign a9980 = a9978 & ~a9632;
assign a9982 = ~a9980 & ~a9626;
assign a9984 = a9982 & ~a9622;
assign a9986 = a9984 & ~a9618;
assign a9988 = a9986 & ~a9614;
assign a9990 = a9988 & ~a9610;
assign a9992 = a9990 & ~a9606;
assign a9994 = a9992 & ~a9598;
assign a9996 = a9994 & ~a9590;
assign a9998 = a9996 & ~a9582;
assign a10000 = a9998 & ~a9574;
assign a10002 = a10000 & ~a9570;
assign a10004 = a10002 & ~a9566;
assign a10006 = a10004 & ~a9560;
assign a10008 = a10006 & ~a9552;
assign a10010 = a10008 & ~a9548;
assign a10012 = a10010 & ~a9544;
assign a10014 = a10012 & ~a9540;
assign a10016 = a10014 & ~a9536;
assign a10018 = a10016 & ~a9532;
assign a10020 = a10018 & ~a9528;
assign a10022 = a10020 & ~a9524;
assign a10024 = a10022 & ~a9516;
assign a10026 = a10024 & ~a9508;
assign a10028 = a10026 & ~a9500;
assign a10030 = a10028 & ~a9492;
assign a10032 = a10030 & ~a9488;
assign a10034 = a10032 & ~a9484;
assign a10036 = a10034 & ~a9480;
assign a10038 = a10036 & ~a9472;
assign a10040 = a10038 & ~a9468;
assign a10042 = a10040 & ~a9462;
assign a10044 = a10042 & ~a9456;
assign a10046 = a10044 & ~a9452;
assign a10048 = a10046 & ~a9448;
assign a10050 = a10048 & ~a9442;
assign a10052 = a10050 & ~a9436;
assign a10054 = a10052 & ~a9432;
assign a10056 = a10054 & ~a9428;
assign a10058 = a10056 & ~a9424;
assign a10060 = a10058 & ~a9420;
assign a10062 = a10060 & ~a9416;
assign a10064 = a10062 & ~a9412;
assign a10066 = a10064 & ~a9408;
assign a10068 = a10066 & ~a9400;
assign a10070 = a10068 & ~a9392;
assign a10072 = a10070 & ~a9384;
assign a10074 = a10072 & ~a9376;
assign a10076 = a10074 & ~a9372;
assign a10078 = a10076 & ~a9368;
assign a10080 = a10078 & ~a9364;
assign a10082 = a10080 & ~a9358;
assign a10084 = a10082 & ~a9352;
assign a10086 = a10084 & ~a9344;
assign a10088 = a10086 & ~a9336;
assign a10090 = a10088 & ~a9328;
assign a10092 = a10090 & ~a9320;
assign a10094 = a9302 & ~l198;
assign a10096 = a10094 & i26;
assign a10098 = a9302 & l186;
assign a10100 = a10098 & ~i14;
assign a10102 = ~a10100 & ~a10096;
assign a10104 = a10102 & ~a10092;
assign a10106 = a10104 & ~a9312;
assign a10108 = ~a10106 & ~a9308;
assign a10110 = a10108 & ~a9300;
assign a10112 = a10110 & ~a9292;
assign a10114 = a10112 & ~a9284;
assign a10116 = a10114 & ~a9276;
assign a10118 = a10116 & ~a9268;
assign a10120 = ~a10118 & ~a9260;
assign a10122 = ~a10120 & ~a9256;
assign a10124 = a10122 & ~a9252;
assign a10126 = a10124 & ~a9248;
assign a10128 = a10126 & ~a9238;
assign a10130 = a10128 & ~a9230;
assign a10132 = a10130 & ~a9222;
assign a10134 = a10132 & ~a9214;
assign a10136 = a10134 & ~a9206;
assign a10138 = a9184 & ~l206;
assign a10140 = a10138 & i34;
assign a10142 = a9184 & ~l204;
assign a10144 = a10142 & i32;
assign a10146 = a9184 & ~l202;
assign a10148 = a10146 & i30;
assign a10150 = a9184 & ~l200;
assign a10152 = a10150 & i28;
assign a10154 = a9184 & ~l198;
assign a10156 = a10154 & i26;
assign a10158 = ~a10156 & ~a10152;
assign a10160 = a10158 & ~a10148;
assign a10162 = a10160 & ~a10144;
assign a10164 = a10162 & ~a10140;
assign a10166 = a10164 & ~a10136;
assign a10168 = a10166 & ~a9198;
assign a10170 = ~a10168 & ~a9194;
assign a10172 = a10170 & ~a9190;
assign a10174 = a10172 & ~a9182;
assign a10176 = a10174 & ~a9178;
assign a10178 = a10176 & ~a9174;
assign a10180 = a10178 & ~a9170;
assign a10182 = a10180 & ~a9166;
assign a10184 = ~a10182 & ~a9162;
assign a10186 = ~a10184 & ~a9158;
assign a10188 = a9068 & ~l216;
assign a10190 = a10188 & ~l208;
assign a10192 = a10190 & i36;
assign a10194 = a10192 & ~l198;
assign a10196 = ~a10194 & ~a10186;
assign a10198 = a10196 & ~a9148;
assign a10200 = ~a10198 & ~a9144;
assign a10202 = a10200 & ~a9140;
assign a10204 = a10202 & ~a9136;
assign a10206 = a10204 & ~a9132;
assign a10208 = a10206 & ~a9124;
assign a10210 = a10208 & ~a9116;
assign a10212 = a10210 & ~a9108;
assign a10214 = ~a10212 & ~a9100;
assign a10216 = ~a10214 & ~a9096;
assign a10218 = a10216 & ~a9092;
assign a10220 = a10218 & ~a9084;
assign a10222 = a10220 & ~a9080;
assign a10224 = a10222 & ~a9074;
assign a10226 = a8996 & ~l216;
assign a10228 = a10226 & ~l208;
assign a10230 = a10228 & i36;
assign a10232 = a10230 & ~l198;
assign a10234 = ~a10232 & ~a10224;
assign a10236 = a10234 & ~a9064;
assign a10238 = ~a10236 & ~a9060;
assign a10240 = a10238 & ~a9056;
assign a10242 = a10240 & ~a9052;
assign a10244 = a10242 & ~a9048;
assign a10246 = a10244 & ~a9044;
assign a10248 = a10246 & ~a9036;
assign a10250 = a10248 & ~a9028;
assign a10252 = a10250 & ~a9020;
assign a10254 = ~a10252 & ~a9012;
assign a10256 = ~a10254 & ~a9008;
assign a10258 = a10256 & ~a9002;
assign a10260 = a10258 & ~a8992;
assign a10262 = a10260 & ~a8988;
assign a10264 = a10262 & ~a8984;
assign a10266 = a10264 & ~a8976;
assign a10268 = a10266 & ~a8968;
assign a10270 = a10268 & ~a8960;
assign a10272 = ~a10270 & ~a8952;
assign a10274 = ~a10272 & ~a8948;
assign a10276 = a10274 & ~a8944;
assign a10278 = a10276 & ~a8940;
assign a10280 = a10278 & ~a8936;
assign a10282 = a8844 & ~l212;
assign a10284 = a10282 & i40;
assign a10286 = ~a10284 & ~a10280;
assign a10288 = a10286 & ~a8924;
assign a10290 = ~a10288 & ~a8920;
assign a10292 = a10290 & ~a8916;
assign a10294 = a10292 & ~a8912;
assign a10296 = a10294 & ~a8908;
assign a10298 = a10296 & ~a8900;
assign a10300 = a10298 & ~a8892;
assign a10302 = a10300 & ~a8884;
assign a10304 = ~a10302 & ~a8876;
assign a10306 = ~a10304 & ~a8872;
assign a10308 = a10306 & ~a8868;
assign a10310 = a10308 & ~a8860;
assign a10312 = a10310 & ~a8856;
assign a10314 = a10312 & ~a8850;
assign a10316 = a7862 & l210;
assign a10318 = a10316 & ~i38;
assign a10320 = ~a10318 & ~a10314;
assign a10322 = a10320 & ~a8842;
assign a10324 = ~a10322 & ~a8838;
assign a10326 = a10324 & ~a8834;
assign a10328 = a10326 & ~a8830;
assign a10330 = a10328 & ~a8826;
assign a10332 = a10330 & ~a8818;
assign a10334 = a10332 & ~a8810;
assign a10336 = a10334 & ~a8802;
assign a10338 = ~a10336 & ~a8794;
assign a10340 = ~a10338 & ~a8790;
assign a10342 = a10340 & ~a8786;
assign a10344 = a10342 & ~a8780;
assign a10346 = a6724 & ~l220;
assign a10348 = a10346 & i48;
assign a10350 = a6724 & ~l218;
assign a10352 = a10350 & i46;
assign a10354 = a6724 & ~l212;
assign a10356 = a10354 & i40;
assign a10358 = a6724 & l214;
assign a10360 = a10358 & ~i42;
assign a10362 = a8770 & ~l214;
assign a10364 = a10362 & i42;
assign a10366 = a10364 & ~l228;
assign a10368 = ~a10366 & ~a10360;
assign a10370 = a10368 & ~a10356;
assign a10372 = a10370 & ~a10352;
assign a10374 = a10372 & ~a10348;
assign a10376 = a10374 & ~a10344;
assign a10378 = a10376 & ~a8774;
assign a10380 = ~a10378 & ~a8768;
assign a10382 = a10380 & ~a8764;
assign a10384 = a10382 & ~a8760;
assign a10386 = a10384 & ~a8756;
assign a10388 = a10386 & ~a8748;
assign a10390 = a10388 & ~a8740;
assign a10392 = a10390 & ~a8732;
assign a10394 = ~a10392 & ~a8724;
assign a10396 = ~a10394 & ~a8720;
assign a10398 = a10396 & ~a8716;
assign a10400 = a10398 & ~a8710;
assign a10402 = a8624 & ~l220;
assign a10404 = a10402 & i48;
assign a10406 = a8624 & ~l212;
assign a10408 = a10406 & i40;
assign a10410 = ~a10408 & ~a10404;
assign a10412 = a10410 & ~a10400;
assign a10414 = a10412 & ~a8706;
assign a10416 = ~a10414 & ~a8700;
assign a10418 = a10416 & ~a8696;
assign a10420 = a10418 & ~a8692;
assign a10422 = a10420 & ~a8688;
assign a10424 = a10422 & ~a8680;
assign a10426 = a10424 & ~a8672;
assign a10428 = a10426 & ~a8664;
assign a10430 = ~a10428 & ~a8656;
assign a10432 = ~a10430 & ~a8652;
assign a10434 = a10432 & ~a8648;
assign a10436 = a10434 & ~a8644;
assign a10438 = a10436 & ~a8636;
assign a10440 = a10438 & ~a8630;
assign a10442 = a8548 & ~l220;
assign a10444 = a10442 & i48;
assign a10446 = a8548 & ~l210;
assign a10448 = a10446 & i38;
assign a10450 = a10448 & ~l228;
assign a10452 = a8548 & l210;
assign a10454 = a10452 & ~i38;
assign a10456 = a8548 & ~l212;
assign a10458 = a10456 & i40;
assign a10460 = a8548 & l214;
assign a10462 = a10460 & ~i42;
assign a10464 = a8548 & ~l214;
assign a10466 = a10464 & i42;
assign a10468 = a10466 & ~l228;
assign a10470 = ~a10468 & ~a10462;
assign a10472 = a10470 & ~a10458;
assign a10474 = a10472 & ~a10454;
assign a10476 = a10474 & ~a10450;
assign a10478 = a10476 & ~a10444;
assign a10480 = a10478 & ~a10440;
assign a10482 = a10480 & ~a8622;
assign a10484 = ~a10482 & ~a8616;
assign a10486 = a10484 & ~a8612;
assign a10488 = a10486 & ~a8608;
assign a10490 = a10488 & ~a8604;
assign a10492 = a10490 & ~a8600;
assign a10494 = a10492 & ~a8596;
assign a10496 = a10494 & ~a8588;
assign a10498 = a10496 & ~a8580;
assign a10500 = a10498 & ~a8572;
assign a10502 = ~a10500 & ~a8564;
assign a10504 = ~a10502 & ~l164;
assign a10506 = a10504 & ~a8560;
assign a10508 = a10506 & ~a8556;
assign a10510 = a8370 & l186;
assign a10512 = a10510 & l204;
assign a10514 = a10512 & ~a8094;
assign a10516 = a10514 & l172;
assign a10518 = a10516 & l170;
assign a10520 = a10518 & ~l168;
assign a10522 = a10520 & ~l166;
assign a10524 = a10522 & l164;
assign a10526 = ~a10524 & ~a10508;
assign a10528 = ~a10526 & ~a8546;
assign a10530 = a10528 & ~a8528;
assign a10532 = ~a10530 & ~a8510;
assign a10534 = a10532 & ~a8492;
assign a10536 = a10534 & ~a8474;
assign a10538 = a10536 & ~a8454;
assign a10540 = ~a10538 & ~a8436;
assign a10542 = a10540 & ~a8422;
assign a10544 = a10542 & ~a8402;
assign a10546 = a10544 & ~a8388;
assign a10548 = ~a10546 & ~a8368;
assign a10550 = a10548 & ~a8354;
assign a10552 = a10550 & ~a8340;
assign a10554 = a10552 & ~a8318;
assign a10556 = a10554 & ~a8300;
assign a10558 = a10556 & ~a8284;
assign a10560 = a10558 & ~a8264;
assign a10562 = a10560 & ~a8246;
assign a10564 = a10562 & ~a8226;
assign a10566 = a10564 & ~a8204;
assign a10568 = ~a10566 & ~a8192;
assign a10570 = a10568 & ~a8174;
assign a10572 = a10570 & ~a8158;
assign a10574 = a10572 & ~a8142;
assign a10576 = a10574 & ~a8128;
assign a10578 = a10576 & ~a8114;
assign a10580 = a10578 & ~a8098;
assign a10582 = ~a10580 & ~a8080;
assign a10584 = a10582 & ~a8064;
assign a10586 = a10584 & ~a8048;
assign a10588 = a10586 & ~a8034;
assign a10590 = ~a10588 & ~a8026;
assign a10592 = a10590 & ~a8002;
assign a10594 = a10592 & ~a7996;
assign a10596 = a10594 & ~a7986;
assign a10598 = a10596 & ~a7976;
assign a10600 = a10598 & ~a7974;
assign a10602 = a10600 & ~a7972;
assign a10604 = a10602 & ~a7970;
assign a10606 = a10604 & ~a7964;
assign a10608 = a10606 & ~a7958;
assign a10610 = a10608 & ~a7946;
assign a10612 = a10610 & ~a7936;
assign a10614 = a10612 & ~a7930;
assign a10616 = a10614 & ~a7920;
assign a10618 = ~a10616 & ~a7918;
assign a10620 = a10618 & ~a7912;
assign a10622 = a10620 & ~a7906;
assign a10624 = a10622 & ~a7900;
assign a10626 = a10624 & ~a7894;
assign a10628 = a10626 & ~a7888;
assign a10630 = a10628 & ~a7882;
assign a10632 = a10630 & ~a7878;
assign a10634 = a10632 & ~a7870;
assign a10636 = a10634 & ~i2;
assign a10638 = ~a10634 & i2;
assign a10640 = ~a10638 & ~a10636;
assign a10642 = a7604 & ~i70;
assign a10644 = a10642 & a7940;
assign a10646 = a8024 & l172;
assign a10648 = a10646 & ~l170;
assign a10650 = a10648 & l168;
assign a10652 = a10650 & l166;
assign a10654 = a10652 & ~l164;
assign a10656 = a8096 & l172;
assign a10658 = a10656 & l170;
assign a10660 = a10658 & ~l168;
assign a10662 = a10660 & ~l166;
assign a10664 = a10662 & l164;
assign a10666 = a8202 & l172;
assign a10668 = a10666 & l170;
assign a10670 = a10668 & ~l168;
assign a10672 = a10670 & ~l166;
assign a10674 = a10672 & l164;
assign a10676 = a8550 & l234;
assign a10678 = a10676 & ~i62;
assign a10680 = a8582 & ~i74;
assign a10682 = a10680 & i72;
assign a10684 = a10682 & ~i70;
assign a10686 = a8550 & ~l214;
assign a10688 = a10686 & i42;
assign a10690 = a10688 & ~l228;
assign a10692 = a8550 & l214;
assign a10694 = a10692 & ~i42;
assign a10696 = a8550 & ~l212;
assign a10698 = a10696 & i40;
assign a10700 = a8550 & l210;
assign a10702 = a10700 & ~i38;
assign a10704 = a8550 & ~l210;
assign a10706 = a10704 & i38;
assign a10708 = a10706 & ~l228;
assign a10710 = a8550 & ~l220;
assign a10712 = a10710 & i48;
assign a10714 = a8550 & ~l216;
assign a10716 = a10714 & l208;
assign a10718 = a10716 & ~i36;
assign a10720 = a8626 & l234;
assign a10722 = a10720 & ~i62;
assign a10724 = a8674 & ~i74;
assign a10726 = a10724 & i72;
assign a10728 = a10726 & ~i70;
assign a10730 = a8626 & ~l212;
assign a10732 = a10730 & i40;
assign a10734 = a8626 & ~l220;
assign a10736 = a10734 & i48;
assign a10738 = a8626 & ~l216;
assign a10740 = a10738 & l208;
assign a10742 = a10740 & ~i36;
assign a10744 = a6726 & l234;
assign a10746 = a10744 & ~i62;
assign a10748 = a8734 & ~i74;
assign a10750 = a10748 & i72;
assign a10752 = a10750 & ~i70;
assign a10754 = a6726 & ~l210;
assign a10756 = a10754 & ~l214;
assign a10758 = a10756 & i42;
assign a10760 = a10758 & ~l228;
assign a10762 = a6726 & l214;
assign a10764 = a10762 & ~i42;
assign a10766 = a6726 & ~l212;
assign a10768 = a10766 & i40;
assign a10770 = a6726 & ~l218;
assign a10772 = a10770 & i46;
assign a10774 = a6726 & ~l220;
assign a10776 = a10774 & i48;
assign a10778 = a10754 & i38;
assign a10780 = a10778 & ~l228;
assign a10782 = a8776 & l234;
assign a10784 = a10782 & ~i62;
assign a10786 = a8804 & ~i74;
assign a10788 = a10786 & i72;
assign a10790 = a10788 & ~i70;
assign a10792 = a8776 & l210;
assign a10794 = a10792 & ~i38;
assign a10796 = a8776 & ~l220;
assign a10798 = a10796 & i48;
assign a10800 = a8846 & l234;
assign a10802 = a10800 & ~i62;
assign a10804 = a8886 & ~i74;
assign a10806 = a10804 & i72;
assign a10808 = a10806 & ~i70;
assign a10810 = a8846 & ~l212;
assign a10812 = a10810 & i40;
assign a10814 = a8846 & ~l220;
assign a10816 = a10814 & i48;
assign a10818 = a8932 & l234;
assign a10820 = a10818 & ~i62;
assign a10822 = a8998 & l234;
assign a10824 = a10822 & ~i62;
assign a10826 = a9030 & ~i74;
assign a10828 = a10826 & i72;
assign a10830 = a10828 & ~i70;
assign a10832 = a8998 & ~l216;
assign a10834 = a10832 & ~l208;
assign a10836 = a10834 & i36;
assign a10838 = a10836 & ~l198;
assign a10840 = a8998 & ~l220;
assign a10842 = a10840 & i48;
assign a10844 = a9070 & l234;
assign a10846 = a10844 & ~i62;
assign a10848 = a9118 & ~i74;
assign a10850 = a10848 & i72;
assign a10852 = a10850 & ~i70;
assign a10854 = a9070 & ~l216;
assign a10856 = a10854 & ~l208;
assign a10858 = a10856 & i36;
assign a10860 = a10858 & ~l198;
assign a10862 = a9070 & ~l220;
assign a10864 = a10862 & i48;
assign a10866 = a9154 & l234;
assign a10868 = a10866 & ~i62;
assign a10870 = a9186 & ~l198;
assign a10872 = a10870 & i26;
assign a10874 = a9186 & ~l200;
assign a10876 = a10874 & i28;
assign a10878 = a9186 & ~l202;
assign a10880 = a10878 & i30;
assign a10882 = a9186 & ~l204;
assign a10884 = a10882 & i32;
assign a10886 = a9186 & ~l206;
assign a10888 = a10886 & i34;
assign a10890 = a9186 & ~l196;
assign a10892 = a10890 & i24;
assign a10894 = a9216 & ~i74;
assign a10896 = a10894 & i72;
assign a10898 = a10896 & ~i70;
assign a10900 = a9244 & l240;
assign a10902 = a10900 & ~i68;
assign a10904 = a9278 & ~i74;
assign a10906 = a10904 & i72;
assign a10908 = a10906 & ~i70;
assign a10910 = a9304 & l186;
assign a10912 = a10910 & ~i14;
assign a10914 = a9304 & ~l198;
assign a10916 = a10914 & i26;
assign a10918 = a9304 & ~l240;
assign a10920 = a10918 & i68;
assign a10922 = a9330 & ~i74;
assign a10924 = a10922 & i72;
assign a10926 = a10924 & ~i70;
assign a10928 = a9394 & ~i74;
assign a10930 = a10928 & i72;
assign a10932 = a10930 & ~i70;
assign a10934 = a9510 & ~i74;
assign a10936 = a10934 & i72;
assign a10938 = a10936 & ~i70;
assign a10940 = a9584 & ~i74;
assign a10942 = a10940 & i72;
assign a10944 = a10942 & ~i70;
assign a10946 = a8928 & ~l164;
assign a10948 = a10946 & ~l210;
assign a10950 = a10948 & i38;
assign a10952 = a10950 & ~l228;
assign a10954 = a9664 & ~i74;
assign a10956 = a10954 & i72;
assign a10958 = a10956 & ~i70;
assign a10960 = a8994 & ~l164;
assign a10962 = a10960 & l214;
assign a10964 = a10962 & ~i42;
assign a10966 = a9150 & ~l164;
assign a10968 = a10966 & l234;
assign a10970 = a10968 & ~i62;
assign a10972 = a10642 & ~a7938;
assign a10974 = ~a10972 & a9750;
assign a10976 = a10974 & ~a9742;
assign a10978 = a10976 & ~a9740;
assign a10980 = a10978 & ~a9738;
assign a10982 = a10980 & ~a9736;
assign a10984 = a10982 & ~a9734;
assign a10986 = a10984 & ~a9732;
assign a10988 = a10986 & ~a9730;
assign a10990 = ~a10988 & ~a10970;
assign a10992 = ~a10990 & ~a9722;
assign a10994 = ~a10992 & a9774;
assign a10996 = a9818 & ~i74;
assign a10998 = a10996 & i72;
assign a11000 = a10998 & ~i70;
assign a11002 = ~a11000 & a9874;
assign a11004 = a11002 & ~a9816;
assign a11006 = a11004 & ~a9808;
assign a11008 = a11006 & ~a9800;
assign a11010 = a11008 & ~a9796;
assign a11012 = a11010 & ~a9792;
assign a11014 = a11012 & ~a9788;
assign a11016 = a11014 & ~a9784;
assign a11018 = a11016 & ~a9780;
assign a11020 = a11018 & ~a10994;
assign a11022 = a11020 & ~a9720;
assign a11024 = a10960 & l210;
assign a11026 = a11024 & ~l214;
assign a11028 = a11026 & i42;
assign a11030 = a11028 & ~l228;
assign a11032 = a10960 & ~l220;
assign a11034 = a11032 & i48;
assign a11036 = a11024 & ~i38;
assign a11038 = ~a11036 & ~a11034;
assign a11040 = a11038 & ~a11030;
assign a11042 = a11040 & ~a11022;
assign a11044 = a11042 & a9712;
assign a11046 = a11044 & ~a10964;
assign a11048 = ~a11046 & ~a9706;
assign a11050 = a11048 & ~a9702;
assign a11052 = a11050 & ~a9698;
assign a11054 = a11052 & ~a9694;
assign a11056 = a11054 & ~a9690;
assign a11058 = a11056 & ~a9686;
assign a11060 = a11058 & ~a9678;
assign a11062 = a11060 & ~a10958;
assign a11064 = a11062 & ~a9662;
assign a11066 = a11064 & ~a9654;
assign a11068 = a11066 & ~a9650;
assign a11070 = a11068 & ~a9646;
assign a11072 = a11070 & ~a9640;
assign a11074 = a10946 & ~l220;
assign a11076 = a11074 & i48;
assign a11078 = a10946 & ~l218;
assign a11080 = a11078 & i46;
assign a11082 = a10946 & ~l212;
assign a11084 = a11082 & i40;
assign a11086 = a10946 & l214;
assign a11088 = a11086 & ~i42;
assign a11090 = a10948 & ~l214;
assign a11092 = a11090 & i42;
assign a11094 = a11092 & ~l228;
assign a11096 = ~a11094 & ~a11088;
assign a11098 = a11096 & ~a11084;
assign a11100 = a11098 & ~a11080;
assign a11102 = a11100 & ~a11076;
assign a11104 = a11102 & ~a11072;
assign a11106 = a11104 & ~a10952;
assign a11108 = ~a11106 & l166;
assign a11110 = a11108 & ~a9626;
assign a11112 = a11110 & ~a9622;
assign a11114 = a11112 & ~a9618;
assign a11116 = a11114 & ~a9614;
assign a11118 = a11116 & ~a9610;
assign a11120 = a11118 & ~a9606;
assign a11122 = a11120 & ~a9598;
assign a11124 = a11122 & ~a10944;
assign a11126 = a11124 & ~a9582;
assign a11128 = a11126 & ~a9574;
assign a11130 = a11128 & ~a9570;
assign a11132 = a11130 & ~a9566;
assign a11134 = a11132 & ~a9560;
assign a11136 = a11134 & ~a9552;
assign a11138 = a11136 & ~a9548;
assign a11140 = a11138 & ~a9544;
assign a11142 = a11140 & ~a9540;
assign a11144 = a11142 & ~a9536;
assign a11146 = a11144 & ~a9532;
assign a11148 = a11146 & ~a9528;
assign a11150 = a11148 & ~a9524;
assign a11152 = a11150 & ~a10938;
assign a11154 = a11152 & ~a9508;
assign a11156 = a11154 & ~a9500;
assign a11158 = a11156 & ~a9492;
assign a11160 = a11158 & ~a9488;
assign a11162 = a11160 & ~a9484;
assign a11164 = a11162 & ~a9480;
assign a11166 = a11164 & ~a9472;
assign a11168 = a11166 & ~a9468;
assign a11170 = a11168 & ~a9462;
assign a11172 = a11170 & ~a9456;
assign a11174 = a11172 & ~a9452;
assign a11176 = a11174 & ~a9448;
assign a11178 = a11176 & ~a9442;
assign a11180 = a11178 & ~a9436;
assign a11182 = a11180 & ~a9432;
assign a11184 = a11182 & ~a9428;
assign a11186 = a11184 & ~a9424;
assign a11188 = a11186 & ~a9420;
assign a11190 = a11188 & ~a9416;
assign a11192 = a11190 & ~a9412;
assign a11194 = a11192 & ~a9408;
assign a11196 = a11194 & ~a10932;
assign a11198 = a11196 & ~a9392;
assign a11200 = a11198 & ~a9384;
assign a11202 = a11200 & ~a9376;
assign a11204 = a11202 & ~a9372;
assign a11206 = a11204 & ~a9368;
assign a11208 = a11206 & ~a9364;
assign a11210 = a11208 & ~a9358;
assign a11212 = a11210 & ~a9352;
assign a11214 = a11212 & ~a9344;
assign a11216 = a11214 & ~a10926;
assign a11218 = a11216 & ~a9328;
assign a11220 = a11218 & ~a9320;
assign a11222 = ~a11220 & ~a10920;
assign a11224 = a11222 & ~a10916;
assign a11226 = a11224 & ~a10912;
assign a11228 = ~a11226 & ~a9308;
assign a11230 = a11228 & ~a9300;
assign a11232 = a11230 & ~a9292;
assign a11234 = a11232 & ~a10908;
assign a11236 = a11234 & ~a9276;
assign a11238 = a11236 & ~a9268;
assign a11240 = ~a11238 & ~a10902;
assign a11242 = ~a11240 & ~a9256;
assign a11244 = a11242 & ~a9252;
assign a11246 = a11244 & ~a9248;
assign a11248 = a11246 & ~a9238;
assign a11250 = a11248 & ~a9230;
assign a11252 = a11250 & ~a10898;
assign a11254 = a11252 & ~a9214;
assign a11256 = a11254 & ~a9206;
assign a11258 = ~a11256 & ~a10892;
assign a11260 = a11258 & ~a10888;
assign a11262 = a11260 & ~a10884;
assign a11264 = a11262 & ~a10880;
assign a11266 = a11264 & ~a10876;
assign a11268 = a11266 & ~a10872;
assign a11270 = ~a11268 & ~a9194;
assign a11272 = a11270 & ~a9190;
assign a11274 = a11272 & ~a9182;
assign a11276 = a11274 & ~a9178;
assign a11278 = a11276 & ~a9174;
assign a11280 = a11278 & ~a9170;
assign a11282 = a11280 & ~a9166;
assign a11284 = ~a11282 & ~a10868;
assign a11286 = ~a11284 & ~a9158;
assign a11288 = ~a11286 & ~a10864;
assign a11290 = a11288 & ~a10860;
assign a11292 = ~a11290 & ~a9144;
assign a11294 = a11292 & ~a9140;
assign a11296 = a11294 & ~a9136;
assign a11298 = a11296 & ~a9132;
assign a11300 = a11298 & ~a10852;
assign a11302 = a11300 & ~a9116;
assign a11304 = a11302 & ~a9108;
assign a11306 = ~a11304 & ~a10846;
assign a11308 = ~a11306 & ~a9096;
assign a11310 = a11308 & ~a9092;
assign a11312 = a11310 & ~a9084;
assign a11314 = a11312 & ~a9080;
assign a11316 = a11314 & ~a9074;
assign a11318 = a11316 & ~a10842;
assign a11320 = ~a11318 & ~a10838;
assign a11322 = ~a11320 & ~a9060;
assign a11324 = a11322 & ~a9056;
assign a11326 = a11324 & ~a9052;
assign a11328 = a11326 & ~a9048;
assign a11330 = a11328 & ~a9044;
assign a11332 = a11330 & ~a10830;
assign a11334 = a11332 & ~a9028;
assign a11336 = a11334 & ~a9020;
assign a11338 = ~a11336 & ~a10824;
assign a11340 = ~a11338 & ~a9008;
assign a11342 = a11340 & ~a9002;
assign a11344 = a11342 & ~a8992;
assign a11346 = a11344 & ~a8988;
assign a11348 = a11346 & ~a8984;
assign a11350 = a11348 & ~a8976;
assign a11352 = a11350 & ~a8968;
assign a11354 = a11352 & ~a8960;
assign a11356 = ~a11354 & ~a10820;
assign a11358 = ~a11356 & ~a8948;
assign a11360 = a11358 & ~a8944;
assign a11362 = a11360 & ~a8940;
assign a11364 = a11362 & ~a8936;
assign a11366 = a11364 & ~a10816;
assign a11368 = a11366 & ~a10812;
assign a11370 = a11368 & ~a8920;
assign a11372 = a11370 & ~a8916;
assign a11374 = a11372 & ~a8912;
assign a11376 = a11374 & ~a8908;
assign a11378 = a11376 & ~a8900;
assign a11380 = a11378 & ~a10808;
assign a11382 = a11380 & ~a8884;
assign a11384 = ~a11382 & ~a10802;
assign a11386 = ~a11384 & ~a8872;
assign a11388 = a11386 & ~a8868;
assign a11390 = a11388 & ~a8860;
assign a11392 = a11390 & ~a8856;
assign a11394 = a11392 & ~a8850;
assign a11396 = a11394 & ~a10798;
assign a11398 = a11396 & ~a10794;
assign a11400 = a11398 & ~a8838;
assign a11402 = a11400 & ~a8834;
assign a11404 = a11402 & ~a8830;
assign a11406 = a11404 & ~a8826;
assign a11408 = a11406 & ~a8818;
assign a11410 = a11408 & ~a10790;
assign a11412 = a11410 & ~a8802;
assign a11414 = ~a11412 & ~a10784;
assign a11416 = ~a11414 & ~a8790;
assign a11418 = a11416 & ~a8786;
assign a11420 = a11418 & ~a8780;
assign a11422 = a11420 & ~a10780;
assign a11424 = a11422 & ~a10776;
assign a11426 = a11424 & ~a10772;
assign a11428 = a11426 & ~a10768;
assign a11430 = a11428 & ~a10764;
assign a11432 = a11430 & ~a10760;
assign a11434 = a11432 & ~a8768;
assign a11436 = a11434 & ~a8764;
assign a11438 = a11436 & ~a8760;
assign a11440 = a11438 & ~a8756;
assign a11442 = a11440 & ~a8748;
assign a11444 = a11442 & ~a10752;
assign a11446 = a11444 & ~a8732;
assign a11448 = ~a11446 & ~a10746;
assign a11450 = ~a11448 & ~a8720;
assign a11452 = a11450 & ~a8716;
assign a11454 = a11452 & ~a8710;
assign a11456 = ~a11454 & ~a10742;
assign a11458 = a11456 & ~a10736;
assign a11460 = a11458 & ~a10732;
assign a11462 = ~a11460 & ~a8700;
assign a11464 = a11462 & ~a8696;
assign a11466 = a11464 & ~a8692;
assign a11468 = a11466 & ~a8688;
assign a11470 = a11468 & ~a10728;
assign a11472 = a11470 & ~a8672;
assign a11474 = a11472 & ~a8664;
assign a11476 = ~a11474 & ~a10722;
assign a11478 = ~a11476 & ~a8652;
assign a11480 = a11478 & ~a8648;
assign a11482 = a11480 & ~a8644;
assign a11484 = a11482 & ~a8636;
assign a11486 = a11484 & ~a8630;
assign a11488 = a11486 & ~a10718;
assign a11490 = ~a11488 & ~a10712;
assign a11492 = a11490 & ~a10708;
assign a11494 = a11492 & ~a10702;
assign a11496 = a11494 & ~a10698;
assign a11498 = a11496 & ~a10694;
assign a11500 = a11498 & ~a10690;
assign a11502 = ~a11500 & ~a8616;
assign a11504 = a11502 & ~a8612;
assign a11506 = a11504 & ~a8608;
assign a11508 = a11506 & ~a8604;
assign a11510 = a11508 & ~a8600;
assign a11512 = a11510 & ~a8596;
assign a11514 = a11512 & ~a10684;
assign a11516 = a11514 & ~a8580;
assign a11518 = a11516 & ~a8572;
assign a11520 = ~a11518 & ~a10678;
assign a11522 = ~a11520 & ~a8560;
assign a11524 = a11522 & ~a8556;
assign a11526 = ~a11524 & ~a10524;
assign a11528 = ~a11526 & ~a8546;
assign a11530 = a11528 & ~a8528;
assign a11532 = ~a11530 & ~a8510;
assign a11534 = a11532 & ~a8492;
assign a11536 = a11534 & ~a8474;
assign a11538 = a11536 & ~a8454;
assign a11540 = ~a11538 & ~a8436;
assign a11542 = a11540 & ~a8422;
assign a11544 = a11542 & ~a8402;
assign a11546 = a11544 & ~a8388;
assign a11548 = a11546 & ~a8368;
assign a11550 = a11548 & ~a8354;
assign a11552 = ~a11550 & ~a8340;
assign a11554 = ~a11552 & ~a8318;
assign a11556 = a11554 & ~a8300;
assign a11558 = a11556 & ~a8284;
assign a11560 = a11558 & ~a8264;
assign a11562 = a11560 & ~a8246;
assign a11564 = ~a11562 & ~a8226;
assign a11566 = a11564 & ~a10674;
assign a11568 = ~a11566 & ~a8192;
assign a11570 = a11568 & ~a8174;
assign a11572 = a11570 & ~a8158;
assign a11574 = a11572 & ~a8142;
assign a11576 = a11574 & ~a8128;
assign a11578 = a11576 & ~a8114;
assign a11580 = a11578 & ~a10664;
assign a11582 = a11580 & ~a8080;
assign a11584 = ~a11582 & ~a8064;
assign a11586 = ~a11584 & ~a8048;
assign a11588 = a11586 & ~a8034;
assign a11590 = a11588 & ~a10654;
assign a11592 = a11590 & ~a8002;
assign a11594 = a11592 & ~a7996;
assign a11596 = a11594 & ~a7986;
assign a11598 = a11596 & ~a7976;
assign a11600 = a11598 & ~a7974;
assign a11602 = a11600 & ~a7972;
assign a11604 = a11602 & ~a7970;
assign a11606 = a11604 & ~a7964;
assign a11608 = a11606 & ~a7958;
assign a11610 = a11608 & ~a10644;
assign a11612 = a11610 & ~a7936;
assign a11614 = a11612 & ~a7930;
assign a11616 = a11614 & ~a7920;
assign a11618 = ~a11616 & ~a7918;
assign a11620 = a11618 & ~a7912;
assign a11622 = a11620 & ~a7906;
assign a11624 = a11622 & ~a7900;
assign a11626 = a11624 & ~a7894;
assign a11628 = a11626 & ~a7888;
assign a11630 = a11628 & ~a7882;
assign a11632 = a11630 & ~a7878;
assign a11634 = a11632 & ~a7870;
assign a11636 = ~a11634 & ~i4;
assign a11638 = a11634 & i4;
assign a11640 = ~a11638 & ~a11636;
assign a11642 = a9556 & ~l210;
assign a11644 = a11642 & ~l214;
assign a11646 = a11644 & i42;
assign a11648 = a11646 & ~l228;
assign a11650 = a9556 & l214;
assign a11652 = a11650 & ~i42;
assign a11654 = a9556 & ~l212;
assign a11656 = a11654 & i40;
assign a11658 = a9556 & ~l218;
assign a11660 = a11658 & i46;
assign a11662 = a9556 & ~l220;
assign a11664 = a11662 & i48;
assign a11666 = a11642 & i38;
assign a11668 = a11666 & ~l228;
assign a11670 = a9636 & l210;
assign a11672 = a11670 & ~i38;
assign a11674 = a9636 & ~l220;
assign a11676 = a11674 & i48;
assign a11678 = a11670 & ~l214;
assign a11680 = a11678 & i42;
assign a11682 = a11680 & ~l228;
assign a11684 = a9636 & l214;
assign a11686 = a11684 & ~i42;
assign a11688 = a9184 & l164;
assign a11690 = a11688 & l236;
assign a11692 = a11690 & ~i64;
assign a11694 = a11688 & l216;
assign a11696 = a11694 & ~l226;
assign a11698 = a11696 & i54;
assign a11700 = a11688 & l214;
assign a11702 = a11700 & ~i42;
assign a11704 = a11688 & ~l210;
assign a11706 = a11704 & i38;
assign a11708 = a11706 & l214;
assign a11710 = a11708 & ~l228;
assign a11712 = a11688 & l186;
assign a11714 = a11712 & ~i14;
assign a11716 = a11688 & l234;
assign a11718 = a11716 & ~i62;
assign a11720 = a7858 & ~l166;
assign a11722 = a11720 & l164;
assign a11724 = a11722 & ~l220;
assign a11726 = a11724 & i48;
assign a11728 = a9724 & ~l164;
assign a11730 = l234 & ~i62;
assign a11732 = ~a11730 & ~a9722;
assign a11734 = a11722 & ~l212;
assign a11736 = a11734 & i40;
assign a11738 = a11722 & ~l196;
assign a11740 = a11738 & i24;
assign a11742 = a11722 & ~l206;
assign a11744 = a11742 & i34;
assign a11746 = a11722 & ~l204;
assign a11748 = a11746 & i32;
assign a11750 = a11722 & ~l202;
assign a11752 = a11750 & i30;
assign a11754 = a11722 & ~l200;
assign a11756 = a11754 & i28;
assign a11758 = a11722 & ~a7960;
assign a11760 = a11758 & ~i74;
assign a11762 = a11760 & ~i72;
assign a11764 = a11762 & i70;
assign a11766 = a11722 & ~a7950;
assign a11768 = a11766 & i74;
assign a11770 = a11768 & i72;
assign a11772 = a11770 & ~i70;
assign a11774 = a11722 & ~a7938;
assign a11776 = a11774 & ~i74;
assign a11778 = a11776 & i72;
assign a11780 = a11778 & ~i70;
assign a11782 = a11722 & ~a7924;
assign a11784 = a11782 & ~i74;
assign a11786 = a11784 & ~i72;
assign a11788 = a11786 & ~i70;
assign a11790 = ~a11788 & ~a11780;
assign a11792 = a11790 & ~a11772;
assign a11794 = a11792 & ~a11764;
assign a11796 = a11794 & ~a11756;
assign a11798 = a11796 & ~a11752;
assign a11800 = a11798 & ~a11748;
assign a11802 = a11800 & ~a11744;
assign a11804 = a11802 & ~a11740;
assign a11806 = a11804 & ~a11736;
assign a11808 = a11806 & ~a11732;
assign a11810 = a11808 & a11728;
assign a11812 = a11810 & ~a11726;
assign a11814 = ~a11812 & ~l168;
assign a11816 = a11814 & ~a11718;
assign a11818 = a11816 & ~a11714;
assign a11820 = a11818 & ~a11710;
assign a11822 = a11820 & ~a11702;
assign a11824 = a11822 & ~a11698;
assign a11826 = a11824 & ~a11692;
assign a11828 = a11826 & ~a11686;
assign a11830 = a11828 & ~a11682;
assign a11832 = a11830 & ~a11676;
assign a11834 = a11832 & ~a11672;
assign a11836 = ~a11834 & ~a9706;
assign a11838 = a11836 & ~a9702;
assign a11840 = a11838 & ~a9698;
assign a11842 = a11840 & ~a9694;
assign a11844 = a11842 & ~a9690;
assign a11846 = a11844 & ~a9686;
assign a11848 = a11846 & ~a9678;
assign a11850 = a11848 & ~a10958;
assign a11852 = a11850 & ~a9662;
assign a11854 = ~a11852 & ~a9654;
assign a11856 = a11854 & ~a9650;
assign a11858 = a11856 & ~a9646;
assign a11860 = a11858 & ~a9640;
assign a11862 = a11860 & ~a11668;
assign a11864 = a11862 & ~a11664;
assign a11866 = a11864 & ~a11660;
assign a11868 = a11866 & ~a11656;
assign a11870 = a11868 & ~a11652;
assign a11872 = a11870 & ~a11648;
assign a11874 = ~a11872 & ~a9626;
assign a11876 = a11874 & ~a9622;
assign a11878 = a11876 & ~a9618;
assign a11880 = a11878 & ~a9614;
assign a11882 = a11880 & ~a9610;
assign a11884 = a11882 & ~a9606;
assign a11886 = a11884 & ~a9598;
assign a11888 = a11886 & ~a10944;
assign a11890 = a11888 & ~a9582;
assign a11892 = ~a11890 & ~a9574;
assign a11894 = a11892 & ~a9570;
assign a11896 = a11894 & ~a9566;
assign a11898 = a11896 & ~a9560;
assign a11900 = ~a11898 & ~a9552;
assign a11902 = a11900 & ~a9548;
assign a11904 = a11902 & ~a9544;
assign a11906 = a11904 & ~a9540;
assign a11908 = a11906 & ~a9536;
assign a11910 = a11908 & ~a9532;
assign a11912 = a11910 & ~a9528;
assign a11914 = a11912 & ~a9524;
assign a11916 = a11914 & ~a10938;
assign a11918 = a11916 & ~a9508;
assign a11920 = a11918 & ~a9500;
assign a11922 = ~a11920 & ~a9492;
assign a11924 = a11922 & ~a9488;
assign a11926 = a11924 & ~a9484;
assign a11928 = a11926 & ~a9480;
assign a11930 = a11928 & ~a9472;
assign a11932 = a11930 & ~a9468;
assign a11934 = a11932 & ~a9462;
assign a11936 = ~a11934 & ~a9456;
assign a11938 = a11936 & ~a9452;
assign a11940 = a11938 & ~a9448;
assign a11942 = a11940 & ~a9442;
assign a11944 = a11942 & ~a9436;
assign a11946 = a11944 & ~a9432;
assign a11948 = a11946 & ~a9428;
assign a11950 = a11948 & ~a9424;
assign a11952 = a11950 & ~a9420;
assign a11954 = a11952 & ~a9416;
assign a11956 = a11954 & ~a9412;
assign a11958 = a11956 & ~a9408;
assign a11960 = a11958 & ~a10932;
assign a11962 = a11960 & ~a9392;
assign a11964 = a11962 & ~a9384;
assign a11966 = ~a11964 & ~a9376;
assign a11968 = a11966 & ~a9372;
assign a11970 = a11968 & ~a9368;
assign a11972 = a11970 & ~a9364;
assign a11974 = a11972 & ~a9358;
assign a11976 = ~a11974 & ~a9352;
assign a11978 = a11976 & ~a9344;
assign a11980 = a11978 & ~a10926;
assign a11982 = a11980 & ~a9328;
assign a11984 = a11982 & ~a9320;
assign a11986 = ~a11984 & ~a10920;
assign a11988 = a11986 & ~a10916;
assign a11990 = a11988 & ~a10912;
assign a11992 = a11990 & ~a9308;
assign a11994 = ~a11992 & ~a9300;
assign a11996 = a11994 & ~a9292;
assign a11998 = a11996 & ~a10908;
assign a12000 = a11998 & ~a9276;
assign a12002 = a12000 & ~a9268;
assign a12004 = ~a12002 & ~a10902;
assign a12006 = a12004 & ~a9256;
assign a12008 = a12006 & ~a9252;
assign a12010 = a12008 & ~a9248;
assign a12012 = ~a12010 & ~a9238;
assign a12014 = a12012 & ~a9230;
assign a12016 = a12014 & ~a10898;
assign a12018 = a12016 & ~a9214;
assign a12020 = a12018 & ~a9206;
assign a12022 = ~a12020 & ~a10892;
assign a12024 = a12022 & ~a10888;
assign a12026 = a12024 & ~a10884;
assign a12028 = a12026 & ~a10880;
assign a12030 = a12028 & ~a10876;
assign a12032 = a12030 & ~a10872;
assign a12034 = a12032 & ~a9194;
assign a12036 = a12034 & ~a9190;
assign a12038 = ~a12036 & ~a9182;
assign a12040 = a12038 & ~a9178;
assign a12042 = a12040 & ~a9174;
assign a12044 = a12042 & ~a9170;
assign a12046 = a12044 & ~a9166;
assign a12048 = ~a12046 & ~a10868;
assign a12050 = a12048 & ~a9158;
assign a12052 = ~a12050 & ~a10864;
assign a12054 = ~a12052 & ~a10860;
assign a12056 = ~a12054 & ~a9144;
assign a12058 = a12056 & ~a9140;
assign a12060 = a12058 & ~a9136;
assign a12062 = a12060 & ~a9132;
assign a12064 = a12062 & ~a10852;
assign a12066 = a12064 & ~a9116;
assign a12068 = a12066 & ~a9108;
assign a12070 = ~a12068 & ~a10846;
assign a12072 = a12070 & ~a9096;
assign a12074 = a12072 & ~a9092;
assign a12076 = a12074 & ~a9084;
assign a12078 = a12076 & ~a9080;
assign a12080 = a12078 & ~a9074;
assign a12082 = a12080 & ~a10842;
assign a12084 = ~a12082 & ~a10838;
assign a12086 = a12084 & ~a9060;
assign a12088 = a12086 & ~a9056;
assign a12090 = a12088 & ~a9052;
assign a12092 = a12090 & ~a9048;
assign a12094 = a12092 & ~a9044;
assign a12096 = a12094 & ~a10830;
assign a12098 = a12096 & ~a9028;
assign a12100 = a12098 & ~a9020;
assign a12102 = ~a12100 & ~a10824;
assign a12104 = a12102 & ~a9008;
assign a12106 = a12104 & ~a9002;
assign a12108 = ~a12106 & ~a8992;
assign a12110 = a12108 & ~a8988;
assign a12112 = a12110 & ~a8984;
assign a12114 = a12112 & ~a8976;
assign a12116 = a12114 & ~a8968;
assign a12118 = a12116 & ~a8960;
assign a12120 = ~a12118 & ~a10820;
assign a12122 = a12120 & ~a8948;
assign a12124 = a12122 & ~a8944;
assign a12126 = a12124 & ~a8940;
assign a12128 = a12126 & ~a8936;
assign a12130 = a12128 & ~a10816;
assign a12132 = a12130 & ~a10812;
assign a12134 = ~a12132 & ~a8920;
assign a12136 = a12134 & ~a8916;
assign a12138 = a12136 & ~a8912;
assign a12140 = a12138 & ~a8908;
assign a12142 = a12140 & ~a8900;
assign a12144 = a12142 & ~a10808;
assign a12146 = a12144 & ~a8884;
assign a12148 = ~a12146 & ~a10802;
assign a12150 = a12148 & ~a8872;
assign a12152 = a12150 & ~a8868;
assign a12154 = a12152 & ~a8860;
assign a12156 = a12154 & ~a8856;
assign a12158 = a12156 & ~a8850;
assign a12160 = a12158 & ~a10798;
assign a12162 = ~a12160 & ~a10794;
assign a12164 = a12162 & ~a8838;
assign a12166 = a12164 & ~a8834;
assign a12168 = a12166 & ~a8830;
assign a12170 = a12168 & ~a8826;
assign a12172 = a12170 & ~a8818;
assign a12174 = a12172 & ~a10790;
assign a12176 = a12174 & ~a8802;
assign a12178 = ~a12176 & ~a10784;
assign a12180 = a12178 & ~a8790;
assign a12182 = a12180 & ~a8786;
assign a12184 = a12182 & ~a8780;
assign a12186 = a12184 & ~a10780;
assign a12188 = ~a12186 & ~a10776;
assign a12190 = a12188 & ~a10772;
assign a12192 = a12190 & ~a10768;
assign a12194 = a12192 & ~a10764;
assign a12196 = a12194 & ~a10760;
assign a12198 = a12196 & ~a8768;
assign a12200 = a12198 & ~a8764;
assign a12202 = a12200 & ~a8760;
assign a12204 = a12202 & ~a8756;
assign a12206 = a12204 & ~a8748;
assign a12208 = a12206 & ~a10752;
assign a12210 = a12208 & ~a8732;
assign a12212 = ~a12210 & ~a10746;
assign a12214 = a12212 & ~a8720;
assign a12216 = a12214 & ~a8716;
assign a12218 = a12216 & ~a8710;
assign a12220 = ~a12218 & ~a10742;
assign a12222 = ~a12220 & ~a10736;
assign a12224 = a12222 & ~a10732;
assign a12226 = ~a12224 & ~a8700;
assign a12228 = a12226 & ~a8696;
assign a12230 = a12228 & ~a8692;
assign a12232 = a12230 & ~a8688;
assign a12234 = a12232 & ~a10728;
assign a12236 = a12234 & ~a8672;
assign a12238 = a12236 & ~a8664;
assign a12240 = ~a12238 & ~a10722;
assign a12242 = a12240 & ~a8652;
assign a12244 = a12242 & ~a8648;
assign a12246 = a12244 & ~a8644;
assign a12248 = a12246 & ~a8636;
assign a12250 = a12248 & ~a8630;
assign a12252 = a12250 & ~a10718;
assign a12254 = ~a12252 & ~a10712;
assign a12256 = a12254 & ~a10708;
assign a12258 = a12256 & ~a10702;
assign a12260 = a12258 & ~a10698;
assign a12262 = a12260 & ~a10694;
assign a12264 = a12262 & ~a10690;
assign a12266 = a12264 & ~a8616;
assign a12268 = a12266 & ~a8612;
assign a12270 = a12268 & ~a8608;
assign a12272 = a12270 & ~a8604;
assign a12274 = a12272 & ~a8600;
assign a12276 = a12274 & ~a8596;
assign a12278 = a12276 & ~a10684;
assign a12280 = a12278 & ~a8580;
assign a12282 = a12280 & ~a8572;
assign a12284 = ~a12282 & ~a10678;
assign a12286 = a12284 & ~a8560;
assign a12288 = a12286 & ~a8556;
assign a12290 = ~a12288 & ~a10524;
assign a12292 = a12290 & ~a8546;
assign a12294 = a12292 & ~a8528;
assign a12296 = ~a12294 & ~a8510;
assign a12298 = a12296 & ~a8492;
assign a12300 = a12298 & ~a8474;
assign a12302 = a12300 & ~a8454;
assign a12304 = ~a12302 & ~a8436;
assign a12306 = a12304 & ~a8422;
assign a12308 = a12306 & ~a8402;
assign a12310 = a12308 & ~a8388;
assign a12312 = a12310 & ~a8368;
assign a12314 = a12312 & ~a8354;
assign a12316 = a12314 & ~a8340;
assign a12318 = ~a12316 & ~a8318;
assign a12320 = a12318 & ~a8300;
assign a12322 = a12320 & ~a8284;
assign a12324 = a12322 & ~a8264;
assign a12326 = ~a12324 & ~a8246;
assign a12328 = ~a12326 & ~a8226;
assign a12330 = ~a12328 & ~a8204;
assign a12332 = ~a12330 & ~a8192;
assign a12334 = a12332 & ~a8174;
assign a12336 = a12334 & ~a8158;
assign a12338 = a12336 & ~a8142;
assign a12340 = a12338 & ~a8128;
assign a12342 = a12340 & ~a8114;
assign a12344 = a12342 & ~a8098;
assign a12346 = ~a12344 & ~a8080;
assign a12348 = a12346 & ~a8064;
assign a12350 = a12348 & ~a8048;
assign a12352 = a12350 & ~a8034;
assign a12354 = ~a12352 & ~a8026;
assign a12356 = ~a12354 & ~a8002;
assign a12358 = a12356 & ~a7996;
assign a12360 = a12358 & ~a7986;
assign a12362 = a12360 & ~a7976;
assign a12364 = a12362 & ~a7974;
assign a12366 = a12364 & ~a7972;
assign a12368 = a12366 & ~a7970;
assign a12370 = a12368 & ~a7964;
assign a12372 = a12370 & ~a7958;
assign a12374 = a12372 & ~a10644;
assign a12376 = a12374 & ~a7936;
assign a12378 = a12376 & ~a7930;
assign a12380 = a12378 & ~a7920;
assign a12382 = ~a12380 & ~a7918;
assign a12384 = a12382 & ~a7912;
assign a12386 = a12384 & ~a7906;
assign a12388 = a12386 & ~a7900;
assign a12390 = a12388 & ~a7894;
assign a12392 = a12390 & ~a7888;
assign a12394 = a12392 & ~a7882;
assign a12396 = a12394 & ~a7878;
assign a12398 = a12396 & ~a7870;
assign a12400 = ~a12398 & ~i6;
assign a12402 = a12398 & i6;
assign a12404 = ~a12402 & ~a12400;
assign a12406 = a11688 & ~a7924;
assign a12408 = a12406 & ~i74;
assign a12410 = a12408 & ~i72;
assign a12412 = a12410 & ~i70;
assign a12414 = a11688 & ~a7938;
assign a12416 = a12414 & ~i70;
assign a12418 = a12416 & ~i74;
assign a12420 = a12418 & i72;
assign a12422 = a11688 & ~a7950;
assign a12424 = a12422 & i74;
assign a12426 = a12424 & i72;
assign a12428 = a12426 & ~i70;
assign a12430 = a11688 & ~a7960;
assign a12432 = a12430 & ~i74;
assign a12434 = a12432 & ~i72;
assign a12436 = a12434 & i70;
assign a12438 = a11688 & ~l200;
assign a12440 = a12438 & i28;
assign a12442 = a11688 & ~l202;
assign a12444 = a12442 & i30;
assign a12446 = a11688 & ~l204;
assign a12448 = a12446 & i32;
assign a12450 = a11688 & ~l206;
assign a12452 = a12450 & i34;
assign a12454 = a11688 & ~l196;
assign a12456 = a12454 & i24;
assign a12458 = a11688 & ~l212;
assign a12460 = a12458 & i40;
assign a12462 = a11688 & ~l220;
assign a12464 = a12462 & i48;
assign a12466 = a11728 & l236;
assign a12468 = a12466 & ~i64;
assign a12470 = a11728 & l234;
assign a12472 = a12470 & ~i62;
assign a12474 = ~a12472 & l170;
assign a12476 = a12474 & ~a12468;
assign a12478 = a12476 & ~a12464;
assign a12480 = a12478 & ~a12460;
assign a12482 = ~a12480 & ~a12456;
assign a12484 = a12482 & ~a12452;
assign a12486 = a12484 & ~a12448;
assign a12488 = a12486 & ~a12444;
assign a12490 = a12488 & ~a12440;
assign a12492 = a12490 & ~a12436;
assign a12494 = a12492 & ~a12428;
assign a12496 = a12494 & ~a12420;
assign a12498 = a12496 & ~a12412;
assign a12500 = ~a12498 & ~a11718;
assign a12502 = a12500 & ~a11714;
assign a12504 = a12502 & ~a11710;
assign a12506 = a12504 & ~a11702;
assign a12508 = a12506 & ~a11698;
assign a12510 = a12508 & ~a11692;
assign a12512 = ~a12510 & ~a11686;
assign a12514 = a12512 & ~a11682;
assign a12516 = a12514 & ~a11676;
assign a12518 = a12516 & ~a11672;
assign a12520 = a12518 & ~a9706;
assign a12522 = a12520 & ~a9702;
assign a12524 = a12522 & ~a9698;
assign a12526 = a12524 & ~a9694;
assign a12528 = a12526 & ~a9690;
assign a12530 = a12528 & ~a9686;
assign a12532 = a12530 & ~a9678;
assign a12534 = a12532 & ~a9670;
assign a12536 = a12534 & ~a9662;
assign a12538 = ~a12536 & ~a9654;
assign a12540 = a12538 & ~a9650;
assign a12542 = a12540 & ~a9646;
assign a12544 = a12542 & ~a9640;
assign a12546 = ~a12544 & ~a11668;
assign a12548 = a12546 & ~a11664;
assign a12550 = a12548 & ~a11660;
assign a12552 = a12550 & ~a11656;
assign a12554 = a12552 & ~a11652;
assign a12556 = a12554 & ~a11648;
assign a12558 = a12556 & ~a9626;
assign a12560 = a12558 & ~a9622;
assign a12562 = a12560 & ~a9618;
assign a12564 = a12562 & ~a9614;
assign a12566 = a12564 & ~a9610;
assign a12568 = a12566 & ~a9606;
assign a12570 = a12568 & ~a9598;
assign a12572 = a12570 & ~a9590;
assign a12574 = a12572 & ~a9582;
assign a12576 = ~a12574 & ~a9574;
assign a12578 = a12576 & ~a9570;
assign a12580 = a12578 & ~a9566;
assign a12582 = a12580 & ~a9560;
assign a12584 = ~a12582 & ~a9552;
assign a12586 = a12584 & ~a9548;
assign a12588 = a12586 & ~a9544;
assign a12590 = a12588 & ~a9540;
assign a12592 = a12590 & ~a9536;
assign a12594 = a12592 & ~a9532;
assign a12596 = a12594 & ~a9528;
assign a12598 = a12596 & ~a9524;
assign a12600 = a12598 & ~a9516;
assign a12602 = a12600 & ~a9508;
assign a12604 = a12602 & ~a9500;
assign a12606 = ~a12604 & ~a9492;
assign a12608 = a12606 & ~a9488;
assign a12610 = a12608 & ~a9484;
assign a12612 = a12610 & ~a9480;
assign a12614 = a12612 & ~a9472;
assign a12616 = a12614 & ~a9468;
assign a12618 = a12616 & ~a9462;
assign a12620 = a12618 & ~a9456;
assign a12622 = a12620 & ~a9452;
assign a12624 = a12622 & ~a9448;
assign a12626 = a12624 & ~a9442;
assign a12628 = a12626 & ~a9436;
assign a12630 = a12628 & ~a9432;
assign a12632 = ~a12630 & ~a9428;
assign a12634 = a12632 & ~a9424;
assign a12636 = a12634 & ~a9420;
assign a12638 = a12636 & ~a9416;
assign a12640 = a12638 & ~a9412;
assign a12642 = a12640 & ~a9408;
assign a12644 = a12642 & ~a9400;
assign a12646 = a12644 & ~a9392;
assign a12648 = a12646 & ~a9384;
assign a12650 = ~a12648 & ~a9376;
assign a12652 = a12650 & ~a9372;
assign a12654 = a12652 & ~a9368;
assign a12656 = a12654 & ~a9364;
assign a12658 = a12656 & ~a9358;
assign a12660 = ~a12658 & ~a9352;
assign a12662 = a12660 & ~a9344;
assign a12664 = a12662 & ~a9336;
assign a12666 = a12664 & ~a9328;
assign a12668 = a12666 & ~a9320;
assign a12670 = ~a12668 & ~a10920;
assign a12672 = a12670 & ~a10916;
assign a12674 = a12672 & ~a10912;
assign a12676 = a12674 & ~a9308;
assign a12678 = ~a12676 & ~a9300;
assign a12680 = a12678 & ~a9292;
assign a12682 = a12680 & ~a9284;
assign a12684 = a12682 & ~a9276;
assign a12686 = a12684 & ~a9268;
assign a12688 = ~a12686 & ~a10902;
assign a12690 = a12688 & ~a9256;
assign a12692 = a12690 & ~a9252;
assign a12694 = a12692 & ~a9248;
assign a12696 = ~a12694 & ~a9238;
assign a12698 = a12696 & ~a9230;
assign a12700 = a12698 & ~a9222;
assign a12702 = a12700 & ~a9214;
assign a12704 = a12702 & ~a9206;
assign a12706 = ~a12704 & ~a10892;
assign a12708 = a12706 & ~a10888;
assign a12710 = a12708 & ~a10884;
assign a12712 = a12710 & ~a10880;
assign a12714 = a12712 & ~a10876;
assign a12716 = a12714 & ~a10872;
assign a12718 = a12716 & ~a9194;
assign a12720 = a12718 & ~a9190;
assign a12722 = ~a12720 & ~a9182;
assign a12724 = a12722 & ~a9178;
assign a12726 = a12724 & ~a9174;
assign a12728 = a12726 & ~a9170;
assign a12730 = a12728 & ~a9166;
assign a12732 = ~a12730 & ~a10868;
assign a12734 = a12732 & ~a9158;
assign a12736 = a12734 & ~a10864;
assign a12738 = a12736 & ~a10860;
assign a12740 = ~a12738 & ~a9144;
assign a12742 = a12740 & ~a9140;
assign a12744 = a12742 & ~a9136;
assign a12746 = a12744 & ~a9132;
assign a12748 = a12746 & ~a9124;
assign a12750 = a12748 & ~a9116;
assign a12752 = a12750 & ~a9108;
assign a12754 = ~a12752 & ~a10846;
assign a12756 = a12754 & ~a9096;
assign a12758 = a12756 & ~a9092;
assign a12760 = a12758 & ~a9084;
assign a12762 = a12760 & ~a9080;
assign a12764 = a12762 & ~a9074;
assign a12766 = ~a12764 & ~a10842;
assign a12768 = a12766 & ~a10838;
assign a12770 = a12768 & ~a9060;
assign a12772 = a12770 & ~a9056;
assign a12774 = a12772 & ~a9052;
assign a12776 = a12774 & ~a9048;
assign a12778 = a12776 & ~a9044;
assign a12780 = a12778 & ~a9036;
assign a12782 = a12780 & ~a9028;
assign a12784 = a12782 & ~a9020;
assign a12786 = ~a12784 & ~a10824;
assign a12788 = a12786 & ~a9008;
assign a12790 = a12788 & ~a9002;
assign a12792 = ~a12790 & ~a8992;
assign a12794 = a12792 & ~a8988;
assign a12796 = a12794 & ~a8984;
assign a12798 = a12796 & ~a8976;
assign a12800 = a12798 & ~a8968;
assign a12802 = a12800 & ~a8960;
assign a12804 = ~a12802 & ~a10820;
assign a12806 = a12804 & ~a8948;
assign a12808 = a12806 & ~a8944;
assign a12810 = a12808 & ~a8940;
assign a12812 = a12810 & ~a8936;
assign a12814 = a12812 & ~a10816;
assign a12816 = a12814 & ~a10812;
assign a12818 = ~a12816 & ~a8920;
assign a12820 = a12818 & ~a8916;
assign a12822 = a12820 & ~a8912;
assign a12824 = a12822 & ~a8908;
assign a12826 = a12824 & ~a8900;
assign a12828 = a12826 & ~a8892;
assign a12830 = a12828 & ~a8884;
assign a12832 = ~a12830 & ~a10802;
assign a12834 = a12832 & ~a8872;
assign a12836 = a12834 & ~a8868;
assign a12838 = a12836 & ~a8860;
assign a12840 = a12838 & ~a8856;
assign a12842 = a12840 & ~a8850;
assign a12844 = a12842 & ~a10798;
assign a12846 = ~a12844 & ~a10794;
assign a12848 = a12846 & ~a8838;
assign a12850 = a12848 & ~a8834;
assign a12852 = a12850 & ~a8830;
assign a12854 = a12852 & ~a8826;
assign a12856 = a12854 & ~a8818;
assign a12858 = a12856 & ~a8810;
assign a12860 = a12858 & ~a8802;
assign a12862 = ~a12860 & ~a10784;
assign a12864 = a12862 & ~a8790;
assign a12866 = a12864 & ~a8786;
assign a12868 = a12866 & ~a8780;
assign a12870 = a12868 & ~a10780;
assign a12872 = ~a12870 & ~a10776;
assign a12874 = a12872 & ~a10772;
assign a12876 = a12874 & ~a10768;
assign a12878 = a12876 & ~a10764;
assign a12880 = a12878 & ~a10760;
assign a12882 = a12880 & ~a8768;
assign a12884 = a12882 & ~a8764;
assign a12886 = a12884 & ~a8760;
assign a12888 = a12886 & ~a8756;
assign a12890 = a12888 & ~a8748;
assign a12892 = a12890 & ~a8740;
assign a12894 = a12892 & ~a8732;
assign a12896 = ~a12894 & ~a10746;
assign a12898 = a12896 & ~a8720;
assign a12900 = a12898 & ~a8716;
assign a12902 = a12900 & ~a8710;
assign a12904 = a12902 & ~a10742;
assign a12906 = a12904 & ~a10736;
assign a12908 = a12906 & ~a10732;
assign a12910 = ~a12908 & ~a8700;
assign a12912 = a12910 & ~a8696;
assign a12914 = a12912 & ~a8692;
assign a12916 = a12914 & ~a8688;
assign a12918 = a12916 & ~a8680;
assign a12920 = a12918 & ~a8672;
assign a12922 = a12920 & ~a8664;
assign a12924 = ~a12922 & ~a10722;
assign a12926 = a12924 & ~a8652;
assign a12928 = a12926 & ~a8648;
assign a12930 = a12928 & ~a8644;
assign a12932 = a12930 & ~a8636;
assign a12934 = a12932 & ~a8630;
assign a12936 = ~a12934 & ~a10718;
assign a12938 = a12936 & ~a10712;
assign a12940 = a12938 & ~a10708;
assign a12942 = a12940 & ~a10702;
assign a12944 = a12942 & ~a10698;
assign a12946 = a12944 & ~a10694;
assign a12948 = a12946 & ~a10690;
assign a12950 = a12948 & ~a8616;
assign a12952 = a12950 & ~a8612;
assign a12954 = a12952 & ~a8608;
assign a12956 = a12954 & ~a8604;
assign a12958 = a12956 & ~a8600;
assign a12960 = a12958 & ~a8596;
assign a12962 = a12960 & ~a8588;
assign a12964 = a12962 & ~a8580;
assign a12966 = a12964 & ~a8572;
assign a12968 = ~a12966 & ~a10678;
assign a12970 = a12968 & ~a8560;
assign a12972 = a12970 & ~a8556;
assign a12974 = ~a12972 & ~a10524;
assign a12976 = ~a12974 & ~a8546;
assign a12978 = a12976 & ~a8528;
assign a12980 = ~a12978 & ~a8510;
assign a12982 = a12980 & ~a8492;
assign a12984 = a12982 & ~a8474;
assign a12986 = a12984 & ~a8454;
assign a12988 = a12986 & ~a8436;
assign a12990 = a12988 & ~a8422;
assign a12992 = ~a12990 & ~a8402;
assign a12994 = a12992 & ~a8388;
assign a12996 = ~a12994 & ~a8368;
assign a12998 = a12996 & ~a8354;
assign a13000 = ~a12998 & ~a8340;
assign a13002 = ~a13000 & ~a8318;
assign a13004 = a13002 & ~a8300;
assign a13006 = ~a13004 & ~a8284;
assign a13008 = a13006 & ~a8264;
assign a13010 = ~a13008 & ~a8246;
assign a13012 = ~a13010 & ~a8226;
assign a13014 = ~a13012 & ~a10674;
assign a13016 = ~a13014 & ~a8192;
assign a13018 = a13016 & ~a8174;
assign a13020 = a13018 & ~a8158;
assign a13022 = a13020 & ~a8142;
assign a13024 = a13022 & ~a8128;
assign a13026 = a13024 & ~a8114;
assign a13028 = a13026 & ~a10664;
assign a13030 = a13028 & ~a8080;
assign a13032 = a13030 & ~a8064;
assign a13034 = a13032 & ~a8048;
assign a13036 = a13034 & ~a8034;
assign a13038 = a13036 & ~a10654;
assign a13040 = ~a13038 & ~a8002;
assign a13042 = a13040 & ~a7996;
assign a13044 = a13042 & ~a7986;
assign a13046 = a13044 & ~a7976;
assign a13048 = a13046 & ~a7974;
assign a13050 = a13048 & ~a7972;
assign a13052 = a13050 & ~a7970;
assign a13054 = a13052 & ~a7964;
assign a13056 = a13054 & ~a7958;
assign a13058 = a13056 & ~a7946;
assign a13060 = a13058 & ~a7936;
assign a13062 = a13060 & ~a7930;
assign a13064 = a13062 & ~a7920;
assign a13066 = ~a13064 & ~a7918;
assign a13068 = a13066 & ~a7912;
assign a13070 = a13068 & ~a7906;
assign a13072 = a13070 & ~a7900;
assign a13074 = a13072 & ~a7894;
assign a13076 = a13074 & ~a7888;
assign a13078 = a13076 & ~a7882;
assign a13080 = a13078 & ~a7878;
assign a13082 = a13080 & ~a7870;
assign a13084 = a13082 & ~i8;
assign a13086 = ~a13082 & i8;
assign a13088 = ~a13086 & ~a13084;
assign a13090 = ~l170 & ~l168;
assign a13092 = a13090 & ~l166;
assign a13094 = a13092 & l164;
assign a13096 = a13094 & l234;
assign a13098 = a13096 & ~i62;
assign a13100 = a13094 & ~l212;
assign a13102 = a13100 & i40;
assign a13104 = a13094 & ~l220;
assign a13106 = a13104 & i48;
assign a13108 = l170 & ~l168;
assign a13110 = a13108 & l166;
assign a13112 = a13110 & ~l164;
assign a13114 = a13112 & l236;
assign a13116 = a13114 & ~i64;
assign a13118 = ~a11730 & ~a9748;
assign a13120 = a13118 & ~a9746;
assign a13122 = a13120 & ~a9744;
assign a13124 = a13122 & ~a9742;
assign a13126 = a13124 & ~a9740;
assign a13128 = a13126 & ~a9738;
assign a13130 = a13128 & ~a9736;
assign a13132 = a13130 & ~a9734;
assign a13134 = a13132 & ~a9732;
assign a13136 = a13134 & ~a9730;
assign a13138 = ~a13136 & a9774;
assign a13140 = a13138 & ~a13116;
assign a13142 = a13140 & ~a13106;
assign a13144 = a13142 & ~a13102;
assign a13146 = ~a13144 & ~a9784;
assign a13148 = a13146 & ~a9788;
assign a13150 = a13148 & ~a9792;
assign a13152 = a13150 & ~a9796;
assign a13154 = a13152 & ~a9800;
assign a13156 = a13154 & ~a9808;
assign a13158 = a13156 & ~a9816;
assign a13160 = a13158 & ~a9824;
assign a13162 = a13160 & ~a9832;
assign a13164 = a13094 & l186;
assign a13166 = a13164 & ~i14;
assign a13168 = a13094 & ~l210;
assign a13170 = a13168 & i38;
assign a13172 = a13170 & l214;
assign a13174 = a13172 & ~l228;
assign a13176 = a13094 & l214;
assign a13178 = a13176 & ~i42;
assign a13180 = a13094 & l216;
assign a13182 = a13180 & ~l226;
assign a13184 = a13182 & i54;
assign a13186 = a13094 & l236;
assign a13188 = a13186 & ~i64;
assign a13190 = ~a13188 & ~a13184;
assign a13192 = a13190 & ~a13178;
assign a13194 = a13192 & ~a13174;
assign a13196 = a13194 & ~a13166;
assign a13198 = a13196 & ~a13162;
assign a13200 = a13198 & a9712;
assign a13202 = a13200 & ~a13098;
assign a13204 = ~a13202 & ~l172;
assign a13206 = a13204 & ~a11686;
assign a13208 = a13206 & ~a11682;
assign a13210 = a13208 & ~a11676;
assign a13212 = ~a13210 & ~a11672;
assign a13214 = ~a13212 & ~a9706;
assign a13216 = a13214 & ~a9702;
assign a13218 = a13216 & ~a9698;
assign a13220 = a13218 & ~a9694;
assign a13222 = a13220 & ~a9690;
assign a13224 = a13222 & ~a9686;
assign a13226 = a13224 & ~a9678;
assign a13228 = a13226 & ~a9670;
assign a13230 = a13228 & ~a9662;
assign a13232 = ~a13230 & ~a9654;
assign a13234 = a13232 & ~a9650;
assign a13236 = a13234 & ~a9646;
assign a13238 = a13236 & ~a9640;
assign a13240 = ~a13238 & ~a11668;
assign a13242 = ~a13240 & ~a11664;
assign a13244 = a13242 & ~a11660;
assign a13246 = a13244 & ~a11656;
assign a13248 = a13246 & ~a11652;
assign a13250 = a13248 & ~a11648;
assign a13252 = ~a13250 & ~a9626;
assign a13254 = a13252 & ~a9622;
assign a13256 = a13254 & ~a9618;
assign a13258 = a13256 & ~a9614;
assign a13260 = a13258 & ~a9610;
assign a13262 = a13260 & ~a9606;
assign a13264 = a13262 & ~a9598;
assign a13266 = a13264 & ~a9590;
assign a13268 = a13266 & ~a9582;
assign a13270 = ~a13268 & ~a9574;
assign a13272 = a13270 & ~a9570;
assign a13274 = a13272 & ~a9566;
assign a13276 = a13274 & ~a9560;
assign a13278 = a13276 & ~a9552;
assign a13280 = a13278 & ~a9548;
assign a13282 = ~a13280 & ~a9544;
assign a13284 = a13282 & ~a9540;
assign a13286 = a13284 & ~a9536;
assign a13288 = a13286 & ~a9532;
assign a13290 = a13288 & ~a9528;
assign a13292 = a13290 & ~a9524;
assign a13294 = a13292 & ~a9516;
assign a13296 = a13294 & ~a9508;
assign a13298 = a13296 & ~a9500;
assign a13300 = ~a13298 & ~a9492;
assign a13302 = a13300 & ~a9488;
assign a13304 = a13302 & ~a9484;
assign a13306 = a13304 & ~a9480;
assign a13308 = a13306 & ~a9472;
assign a13310 = a13308 & ~a9468;
assign a13312 = a13310 & ~a9462;
assign a13314 = ~a13312 & ~a9456;
assign a13316 = a13314 & ~a9452;
assign a13318 = a13316 & ~a9448;
assign a13320 = a13318 & ~a9442;
assign a13322 = a13320 & ~a9436;
assign a13324 = a13322 & ~a9432;
assign a13326 = a13324 & ~a9428;
assign a13328 = a13326 & ~a9424;
assign a13330 = a13328 & ~a9420;
assign a13332 = a13330 & ~a9416;
assign a13334 = a13332 & ~a9412;
assign a13336 = a13334 & ~a9408;
assign a13338 = a13336 & ~a9400;
assign a13340 = a13338 & ~a9392;
assign a13342 = a13340 & ~a9384;
assign a13344 = ~a13342 & ~a9376;
assign a13346 = a13344 & ~a9372;
assign a13348 = a13346 & ~a9368;
assign a13350 = a13348 & ~a9364;
assign a13352 = a13350 & ~a9358;
assign a13354 = ~a13352 & ~a9352;
assign a13356 = a13354 & ~a9344;
assign a13358 = a13356 & ~a9336;
assign a13360 = a13358 & ~a9328;
assign a13362 = a13360 & ~a9320;
assign a13364 = a13362 & ~a10920;
assign a13366 = a13364 & ~a10916;
assign a13368 = a13366 & ~a10912;
assign a13370 = ~a13368 & ~a9308;
assign a13372 = ~a13370 & ~a9300;
assign a13374 = a13372 & ~a9292;
assign a13376 = a13374 & ~a9284;
assign a13378 = a13376 & ~a9276;
assign a13380 = a13378 & ~a9268;
assign a13382 = a13380 & ~a10902;
assign a13384 = ~a13382 & ~a9256;
assign a13386 = a13384 & ~a9252;
assign a13388 = a13386 & ~a9248;
assign a13390 = ~a13388 & ~a9238;
assign a13392 = a13390 & ~a9230;
assign a13394 = a13392 & ~a9222;
assign a13396 = a13394 & ~a9214;
assign a13398 = a13396 & ~a9206;
assign a13400 = a13398 & ~a10892;
assign a13402 = a13400 & ~a10888;
assign a13404 = a13402 & ~a10884;
assign a13406 = a13404 & ~a10880;
assign a13408 = a13406 & ~a10876;
assign a13410 = a13408 & ~a10872;
assign a13412 = ~a13410 & ~a9194;
assign a13414 = a13412 & ~a9190;
assign a13416 = ~a13414 & ~a9182;
assign a13418 = a13416 & ~a9178;
assign a13420 = a13418 & ~a9174;
assign a13422 = a13420 & ~a9170;
assign a13424 = a13422 & ~a9166;
assign a13426 = a13424 & ~a10868;
assign a13428 = ~a13426 & ~a9158;
assign a13430 = a13428 & ~a10864;
assign a13432 = a13430 & ~a10860;
assign a13434 = ~a13432 & ~a9144;
assign a13436 = a13434 & ~a9140;
assign a13438 = a13436 & ~a9136;
assign a13440 = a13438 & ~a9132;
assign a13442 = a13440 & ~a9124;
assign a13444 = a13442 & ~a9116;
assign a13446 = a13444 & ~a9108;
assign a13448 = a13446 & ~a10846;
assign a13450 = ~a13448 & ~a9096;
assign a13452 = a13450 & ~a9092;
assign a13454 = a13452 & ~a9084;
assign a13456 = a13454 & ~a9080;
assign a13458 = a13456 & ~a9074;
assign a13460 = ~a13458 & ~a10842;
assign a13462 = a13460 & ~a10838;
assign a13464 = a13462 & ~a9060;
assign a13466 = a13464 & ~a9056;
assign a13468 = a13466 & ~a9052;
assign a13470 = a13468 & ~a9048;
assign a13472 = a13470 & ~a9044;
assign a13474 = a13472 & ~a9036;
assign a13476 = a13474 & ~a9028;
assign a13478 = a13476 & ~a9020;
assign a13480 = a13478 & ~a10824;
assign a13482 = ~a13480 & ~a9008;
assign a13484 = a13482 & ~a9002;
assign a13486 = ~a13484 & ~a8992;
assign a13488 = a13486 & ~a8988;
assign a13490 = a13488 & ~a8984;
assign a13492 = a13490 & ~a8976;
assign a13494 = a13492 & ~a8968;
assign a13496 = a13494 & ~a8960;
assign a13498 = a13496 & ~a10820;
assign a13500 = ~a13498 & ~a8948;
assign a13502 = a13500 & ~a8944;
assign a13504 = a13502 & ~a8940;
assign a13506 = a13504 & ~a8936;
assign a13508 = ~a13506 & ~a10816;
assign a13510 = a13508 & ~a10812;
assign a13512 = a13510 & ~a8920;
assign a13514 = a13512 & ~a8916;
assign a13516 = a13514 & ~a8912;
assign a13518 = a13516 & ~a8908;
assign a13520 = a13518 & ~a8900;
assign a13522 = a13520 & ~a8892;
assign a13524 = a13522 & ~a8884;
assign a13526 = a13524 & ~a10802;
assign a13528 = ~a13526 & ~a8872;
assign a13530 = a13528 & ~a8868;
assign a13532 = a13530 & ~a8860;
assign a13534 = a13532 & ~a8856;
assign a13536 = a13534 & ~a8850;
assign a13538 = a13536 & ~a10798;
assign a13540 = ~a13538 & ~a10794;
assign a13542 = a13540 & ~a8838;
assign a13544 = a13542 & ~a8834;
assign a13546 = a13544 & ~a8830;
assign a13548 = a13546 & ~a8826;
assign a13550 = a13548 & ~a8818;
assign a13552 = a13550 & ~a8810;
assign a13554 = a13552 & ~a8802;
assign a13556 = a13554 & ~a10784;
assign a13558 = ~a13556 & ~a8790;
assign a13560 = a13558 & ~a8786;
assign a13562 = a13560 & ~a8780;
assign a13564 = a13562 & ~a10780;
assign a13566 = ~a13564 & ~a10776;
assign a13568 = a13566 & ~a10772;
assign a13570 = a13568 & ~a10768;
assign a13572 = a13570 & ~a10764;
assign a13574 = a13572 & ~a10760;
assign a13576 = a13574 & ~a8768;
assign a13578 = a13576 & ~a8764;
assign a13580 = a13578 & ~a8760;
assign a13582 = a13580 & ~a8756;
assign a13584 = a13582 & ~a8748;
assign a13586 = a13584 & ~a8740;
assign a13588 = a13586 & ~a8732;
assign a13590 = a13588 & ~a10746;
assign a13592 = ~a13590 & ~a8720;
assign a13594 = a13592 & ~a8716;
assign a13596 = a13594 & ~a8710;
assign a13598 = a13596 & ~a10742;
assign a13600 = a13598 & ~a10736;
assign a13602 = a13600 & ~a10732;
assign a13604 = ~a13602 & ~a8700;
assign a13606 = a13604 & ~a8696;
assign a13608 = a13606 & ~a8692;
assign a13610 = a13608 & ~a8688;
assign a13612 = a13610 & ~a8680;
assign a13614 = a13612 & ~a8672;
assign a13616 = a13614 & ~a8664;
assign a13618 = a13616 & ~a10722;
assign a13620 = ~a13618 & ~a8652;
assign a13622 = a13620 & ~a8648;
assign a13624 = a13622 & ~a8644;
assign a13626 = a13624 & ~a8636;
assign a13628 = a13626 & ~a8630;
assign a13630 = ~a13628 & ~a10718;
assign a13632 = a13630 & ~a10712;
assign a13634 = a13632 & ~a10708;
assign a13636 = a13634 & ~a10702;
assign a13638 = a13636 & ~a10698;
assign a13640 = a13638 & ~a10694;
assign a13642 = a13640 & ~a10690;
assign a13644 = a13642 & ~a8616;
assign a13646 = a13644 & ~a8612;
assign a13648 = a13646 & ~a8608;
assign a13650 = a13648 & ~a8604;
assign a13652 = a13650 & ~a8600;
assign a13654 = a13652 & ~a8596;
assign a13656 = a13654 & ~a8588;
assign a13658 = a13656 & ~a8580;
assign a13660 = a13658 & ~a8572;
assign a13662 = a13660 & ~a10678;
assign a13664 = ~a13662 & ~a8560;
assign a13666 = a13664 & ~a8556;
assign a13668 = a13666 & ~a10524;
assign a13670 = a13668 & ~a8546;
assign a13672 = a13670 & ~a8528;
assign a13674 = ~a13672 & ~a8510;
assign a13676 = a13674 & ~a8492;
assign a13678 = ~a13676 & ~a8474;
assign a13680 = a13678 & ~a8454;
assign a13682 = a13680 & ~a8436;
assign a13684 = a13682 & ~a8422;
assign a13686 = ~a13684 & ~a8402;
assign a13688 = a13686 & ~a8388;
assign a13690 = ~a13688 & ~a8368;
assign a13692 = a13690 & ~a8354;
assign a13694 = a13692 & ~a8340;
assign a13696 = ~a13694 & ~a8318;
assign a13698 = ~a13696 & ~a8300;
assign a13700 = ~a13698 & ~a8284;
assign a13702 = ~a13700 & ~a8264;
assign a13704 = ~a13702 & ~a8246;
assign a13706 = ~a13704 & ~a8226;
assign a13708 = ~a13706 & ~a10674;
assign a13710 = ~a13708 & ~a8192;
assign a13712 = a13710 & ~a8174;
assign a13714 = a13712 & ~a8158;
assign a13716 = a13714 & ~a8142;
assign a13718 = a13716 & ~a8128;
assign a13720 = a13718 & ~a8114;
assign a13722 = a13720 & ~a10664;
assign a13724 = ~a13722 & ~a8080;
assign a13726 = a13724 & ~a8064;
assign a13728 = ~a13726 & ~a8048;
assign a13730 = a13728 & ~a8034;
assign a13732 = a13730 & ~a10654;
assign a13734 = ~a13732 & ~a8002;
assign a13736 = a13734 & ~a7996;
assign a13738 = a13736 & ~a7986;
assign a13740 = a13738 & ~a7976;
assign a13742 = a13740 & ~a7974;
assign a13744 = a13742 & ~a7972;
assign a13746 = a13744 & ~a7970;
assign a13748 = a13746 & ~a7964;
assign a13750 = a13748 & ~a7958;
assign a13752 = a13750 & ~a7946;
assign a13754 = a13752 & ~a7936;
assign a13756 = a13754 & ~a7930;
assign a13758 = a13756 & ~a7920;
assign a13760 = a13758 & ~a7918;
assign a13762 = a13760 & ~a7912;
assign a13764 = a13762 & ~a7906;
assign a13766 = a13764 & ~a7900;
assign a13768 = a13766 & ~a7894;
assign a13770 = a13768 & ~a7888;
assign a13772 = a13770 & ~a7882;
assign a13774 = a13772 & ~a7878;
assign a13776 = a13774 & ~a7870;
assign a13778 = ~a13776 & ~i10;
assign a13780 = a13776 & i10;
assign a13782 = ~a13780 & ~a13778;
assign a13784 = ~i102 & ~i100;
assign a13786 = a13784 & ~a2238;
assign a13788 = i102 & i100;
assign a13790 = a13788 & ~a2306;
assign a13792 = ~a13790 & ~a13786;
assign a13794 = ~a13792 & i104;
assign a13796 = ~i104 & ~i102;
assign a13798 = a13796 & ~i100;
assign a13800 = a13798 & ~a2384;
assign a13802 = ~i104 & i102;
assign a13804 = a13802 & i100;
assign a13806 = a13804 & ~a2520;
assign a13808 = ~a13806 & ~a13800;
assign a13810 = a13808 & ~a13794;
assign a13812 = ~a13810 & i98;
assign a13814 = i104 & ~i102;
assign a13816 = a13814 & i100;
assign a13818 = a13816 & ~i98;
assign a13820 = a13818 & ~a4346;
assign a13822 = ~a13820 & ~a13812;
assign a13824 = ~a13822 & ~i96;
assign a13826 = a13798 & ~i98;
assign a13828 = a13826 & i96;
assign a13830 = a13828 & ~a1450;
assign a13832 = i104 & i102;
assign a13834 = a13832 & ~i100;
assign a13836 = a13834 & i98;
assign a13838 = a13836 & ~i96;
assign a13840 = a13838 & ~a1514;
assign a13842 = a13802 & ~i100;
assign a13844 = a13842 & i98;
assign a13846 = a13844 & ~i96;
assign a13848 = a13846 & ~a1652;
assign a13850 = a13834 & ~i98;
assign a13852 = a13850 & ~i96;
assign a13854 = a13852 & ~a1774;
assign a13856 = a13832 & i100;
assign a13858 = a13856 & ~i98;
assign a13860 = a13858 & ~i96;
assign a13862 = a13860 & ~a1898;
assign a13864 = a13796 & i100;
assign a13866 = a13864 & ~i98;
assign a13868 = a13866 & ~i96;
assign a13870 = a13868 & ~a6030;
assign a13872 = ~l320 & ~l318;
assign a13874 = ~a13872 & ~a13870;
assign a13876 = a13874 & ~a13862;
assign a13878 = a13876 & ~a13854;
assign a13880 = a13878 & ~a13848;
assign a13882 = a13880 & ~a13840;
assign a13884 = a13882 & ~a13830;
assign a13886 = a13884 & ~a13824;
assign a13888 = ~a13886 & i146;
assign a13890 = a13886 & ~i146;
assign a13892 = ~a13890 & ~a13888;
assign a13894 = ~l316 & ~l314;
assign a13896 = ~a13894 & ~a13870;
assign a13898 = a13896 & ~a13862;
assign a13900 = a13898 & ~a13854;
assign a13902 = a13900 & ~a13848;
assign a13904 = a13902 & ~a13840;
assign a13906 = a13904 & ~a13830;
assign a13908 = a13906 & ~a13824;
assign a13910 = ~a13908 & i142;
assign a13912 = a13908 & ~i142;
assign a13914 = ~a13912 & ~a13910;
assign a13916 = l334 & l332;
assign a13918 = a13916 & l336;
assign a13920 = ~a13918 & ~l324;
assign a13922 = ~a13920 & ~a13870;
assign a13924 = a13922 & ~a13862;
assign a13926 = a13924 & ~a13854;
assign a13928 = a13926 & ~a13848;
assign a13930 = a13928 & ~a13840;
assign a13932 = a13930 & ~a13830;
assign a13934 = a13932 & ~a13824;
assign a13936 = ~a13934 & i150;
assign a13938 = a13934 & ~i150;
assign a13940 = ~a13938 & ~a13936;
assign a13942 = ~a13916 & ~l326;
assign a13944 = ~a13942 & ~a13870;
assign a13946 = a13944 & ~a13862;
assign a13948 = a13946 & ~a13854;
assign a13950 = a13948 & ~a13848;
assign a13952 = a13950 & ~a13840;
assign a13954 = a13952 & ~a13830;
assign a13956 = a13954 & ~a13824;
assign a13958 = ~a13956 & i152;
assign a13960 = a13956 & ~i152;
assign a13962 = ~a13960 & ~a13958;
assign a13964 = ~a13792 & i98;
assign a13966 = ~i102 & i100;
assign a13968 = a13966 & ~i98;
assign a13970 = a13968 & ~a4346;
assign a13972 = ~a13970 & ~a13964;
assign a13974 = i104 & ~i96;
assign a13976 = a13974 & ~a13972;
assign a13978 = a13918 & l322;
assign a13980 = ~a13978 & ~l328;
assign a13982 = ~a13980 & ~a13976;
assign a13984 = a13982 & ~a13830;
assign a13986 = a13984 & ~a13840;
assign a13988 = a13986 & ~a13848;
assign a13990 = a13988 & ~a13854;
assign a13992 = a13990 & ~a13862;
assign a13994 = a13992 & ~a13870;
assign a13996 = a13994 & ~i154;
assign a13998 = ~a13994 & i154;
assign a14000 = ~a13998 & ~a13996;
assign a14002 = a13802 & i98;
assign a14004 = a14002 & ~a2520;
assign a14006 = a13814 & ~i98;
assign a14008 = a14006 & ~a4346;
assign a14010 = ~a14008 & ~a14004;
assign a14012 = i100 & ~i96;
assign a14014 = a14012 & ~a14010;
assign a14016 = ~l336 & ~l330;
assign a14018 = ~a14016 & ~a14014;
assign a14020 = a14018 & ~a13830;
assign a14022 = a14020 & ~a13840;
assign a14024 = a14022 & ~a13848;
assign a14026 = a14024 & ~a13854;
assign a14028 = a14026 & ~a13862;
assign a14030 = a14028 & ~a13870;
assign a14032 = a14030 & ~i156;
assign a14034 = ~a14030 & i156;
assign a14036 = ~a14034 & ~a14032;
assign a14038 = ~l236 & i64;
assign a14040 = a14038 & l312;
assign a14042 = l312 & ~i140;
assign a14044 = ~a14042 & l310;
assign a14046 = ~a14044 & ~a14040;
assign a14048 = a14046 & i138;
assign a14050 = ~a14046 & ~i138;
assign a14052 = ~a14050 & ~a14048;
assign a14054 = a13798 & i98;
assign a14056 = a14054 & ~i96;
assign a14058 = ~a14056 & a2384;
assign a14060 = a14056 & ~a2384;
assign a14062 = ~a14060 & l312;
assign a14064 = ~a14062 & ~a14058;
assign a14066 = ~a14064 & ~i140;
assign a14068 = a14064 & i140;
assign a14070 = ~a14068 & ~a14066;
assign a14072 = ~l192 & l190;
assign a14074 = a14072 & l188;
assign a14076 = a14074 & ~l204;
assign a14078 = ~a14074 & l204;
assign a14080 = ~a14078 & ~a14076;
assign a14082 = ~l192 & ~l190;
assign a14084 = a14082 & ~l188;
assign a14086 = a14084 & ~l202;
assign a14088 = ~a14084 & l202;
assign a14090 = ~a14088 & ~a14086;
assign a14092 = l192 & l190;
assign a14094 = a14092 & ~l188;
assign a14096 = a14094 & ~l206;
assign a14098 = ~a14094 & l206;
assign a14100 = ~a14098 & ~a14096;
assign a14102 = a14072 & ~l188;
assign a14104 = a14102 & ~l200;
assign a14106 = ~a14102 & l200;
assign a14108 = ~a14106 & ~a14104;
assign a14110 = a14082 & l188;
assign a14112 = a14110 & ~l198;
assign a14114 = ~a14110 & l198;
assign a14116 = ~a14114 & ~a14112;
assign a14118 = ~a6676 & ~l242;
assign a14120 = ~a14118 & ~a7960;
assign a14122 = a14120 & ~a7932;
assign a14124 = ~a14122 & ~l234;
assign a14126 = a14122 & l234;
assign a14128 = ~a14126 & ~a14124;
assign a14130 = ~l206 & ~l194;
assign a14132 = a14130 & l186;
assign a14134 = a14132 & ~l196;
assign a14136 = ~a14132 & l196;
assign a14138 = ~a14136 & ~a14134;
assign a14140 = l266 & ~l230;
assign a14142 = ~a14140 & a7060;
assign a14144 = a14142 & ~l218;
assign a14146 = ~a14142 & l218;
assign a14148 = ~a14146 & ~a14144;
assign a14150 = l192 & ~l190;
assign a14152 = a14150 & l188;
assign a14154 = ~a14152 & l184;
assign a14156 = a14154 & ~l186;
assign a14158 = ~a14154 & l186;
assign a14160 = ~a14158 & ~a14156;
assign a14162 = ~l204 & ~l198;
assign a14164 = a14162 & ~l200;
assign a14166 = a14164 & ~l202;
assign a14168 = ~a14166 & ~l194;
assign a14170 = a14166 & l194;
assign a14172 = ~a14170 & ~a14168;
assign a14174 = l294 & ~l292;
assign a14176 = ~a14084 & ~l184;
assign a14178 = ~l284 & i112;
assign a14180 = l284 & ~i112;
assign a14182 = ~a14180 & ~a14178;
assign a14184 = ~a14038 & ~a9722;
assign a14186 = ~l286 & i114;
assign a14188 = l286 & ~i114;
assign a14190 = ~a14188 & ~a14186;
assign a14192 = ~l216 & i44;
assign a14194 = l216 & ~i44;
assign a14196 = ~a14194 & ~a14192;
assign a14198 = ~l238 & i66;
assign a14200 = l238 & ~i66;
assign a14202 = ~a14200 & ~a14198;
assign a14204 = ~l288 & i116;
assign a14206 = l288 & ~i116;
assign a14208 = ~a14206 & ~a14204;
assign a14210 = ~l290 & i118;
assign a14212 = l290 & ~i118;
assign a14214 = ~a14212 & ~a14210;
assign a14216 = ~l282 & i110;
assign a14218 = l282 & ~i110;
assign a14220 = ~a14218 & ~a14216;
assign a14222 = ~l280 & i108;
assign a14224 = l280 & ~i108;
assign a14226 = ~a14224 & ~a14222;
assign a14228 = ~l278 & i106;
assign a14230 = l278 & ~i106;
assign a14232 = ~a14230 & ~a14228;
assign a14234 = ~l296 & i124;
assign a14236 = l296 & ~i124;
assign a14238 = ~a14236 & ~a14234;
assign a14240 = l298 & ~i126;
assign a14242 = ~a14240 & ~a3560;
assign a14244 = ~l300 & i128;
assign a14246 = l300 & ~i128;
assign a14248 = ~a14246 & ~a14244;
assign a14250 = ~l294 & i122;
assign a14252 = l294 & ~i122;
assign a14254 = ~a14252 & ~a14250;
assign a14256 = ~l292 & i120;
assign a14258 = l292 & ~i120;
assign a14260 = ~a14258 & ~a14256;
assign a14262 = ~l302 & i130;
assign a14264 = l302 & ~i130;
assign a14266 = ~a14264 & ~a14262;
assign a14268 = ~l304 & i132;
assign a14270 = l304 & ~i132;
assign a14272 = ~a14270 & ~a14268;
assign a14274 = ~l306 & i134;
assign a14276 = l306 & ~i134;
assign a14278 = ~a14276 & ~a14274;
assign a14280 = ~l308 & i136;
assign a14282 = l308 & ~i136;
assign a14284 = ~a14282 & ~a14280;
assign a14286 = ~l260 & i88;
assign a14288 = ~a14286 & ~a7660;
assign a14290 = ~l262 & i90;
assign a14292 = ~a14290 & ~a7658;
assign a14294 = ~l258 & i86;
assign a14296 = l258 & ~i86;
assign a14298 = ~a14296 & ~a14294;
assign a14300 = ~l256 & i84;
assign a14302 = l256 & ~i84;
assign a14304 = ~a14302 & ~a14300;
assign a14306 = ~l254 & i82;
assign a14308 = l254 & ~i82;
assign a14310 = ~a14308 & ~a14306;
assign a14312 = ~l266 & i94;
assign a14314 = l266 & ~i94;
assign a14316 = ~a14314 & ~a14312;
assign a14318 = l264 & ~i92;
assign a14320 = ~a14318 & ~a7652;
assign a14322 = ~l232 & i60;
assign a14324 = l232 & ~i60;
assign a14326 = ~a14324 & ~a14322;
assign a14328 = ~l208 & i36;
assign a14330 = l208 & ~i36;
assign a14332 = ~a14330 & ~a14328;
assign a14334 = l240 & ~i68;
assign a14336 = ~a14334 & ~a7664;
assign a14338 = ~l210 & i38;
assign a14340 = l210 & ~i38;
assign a14342 = ~a14340 & ~a14338;
assign a14344 = ~l212 & i40;
assign a14346 = l212 & ~i40;
assign a14348 = ~a14346 & ~a14344;
assign a14350 = ~l214 & i42;
assign a14352 = l214 & ~i42;
assign a14354 = ~a14352 & ~a14350;
assign a14356 = ~l246 & i74;
assign a14358 = l246 & ~i74;
assign a14360 = ~a14358 & ~a14356;
assign a14362 = ~l244 & i72;
assign a14364 = l244 & ~i72;
assign a14366 = ~a14364 & ~a14362;
assign a14368 = ~l242 & i70;
assign a14370 = l242 & ~i70;
assign a14372 = ~a14370 & ~a14368;
assign a14374 = ~l220 & i48;
assign a14376 = l220 & ~i48;
assign a14378 = ~a14376 & ~a14374;
assign a14380 = ~l222 & i50;
assign a14382 = l222 & ~i50;
assign a14384 = ~a14382 & ~a14380;
assign a14386 = ~l224 & i52;
assign a14388 = l224 & ~i52;
assign a14390 = ~a14388 & ~a14386;
assign a14392 = ~l228 & i56;
assign a14394 = l228 & ~i56;
assign a14396 = ~a14394 & ~a14392;
assign a14398 = ~l226 & i54;
assign a14400 = l226 & ~i54;
assign a14402 = ~a14400 & ~a14398;
assign a14404 = ~l230 & i58;
assign a14406 = l230 & ~i58;
assign a14408 = ~a14406 & ~a14404;
assign a14410 = ~l192 & i20;
assign a14412 = l192 & ~i20;
assign a14414 = ~a14412 & ~a14410;
assign a14416 = ~l190 & i18;
assign a14418 = l190 & ~i18;
assign a14420 = ~a14418 & ~a14416;
assign a14422 = ~l188 & i16;
assign a14424 = l188 & ~i16;
assign a14426 = ~a14424 & ~a14422;
assign a14428 = l184 & ~i12;
assign a14430 = ~a14428 & ~a7662;
assign a14432 = ~l336 & ~i162;
assign a14434 = l336 & i162;
assign a14436 = ~a14434 & ~a14432;
assign a14438 = ~l334 & ~i160;
assign a14440 = l334 & i160;
assign a14442 = ~a14440 & ~a14438;
assign a14444 = ~l334 & i160;
assign a14446 = l334 & ~i160;
assign a14448 = ~a14446 & ~a14444;
assign a14450 = ~l332 & ~i158;
assign a14452 = l332 & i158;
assign a14454 = ~a14452 & ~a14450;
assign a14456 = a14454 & a14448;
assign a14458 = ~a14456 & ~a14442;
assign a14460 = ~a14458 & a14436;
assign a14462 = ~l336 & i162;
assign a14464 = l336 & ~i162;
assign a14466 = ~a14464 & ~a14462;
assign a14468 = a14454 & a14442;
assign a14470 = a14468 & a14466;
assign a14472 = ~a14470 & ~a14460;
assign a14474 = ~a14472 & a14430;
assign a14476 = ~l184 & ~i12;
assign a14478 = l184 & i12;
assign a14480 = ~a14478 & ~a14476;
assign a14482 = ~l332 & i158;
assign a14484 = l332 & ~i158;
assign a14486 = ~a14484 & ~a14482;
assign a14488 = a14486 & a14448;
assign a14490 = a14488 & a14466;
assign a14492 = a14490 & a14480;
assign a14494 = ~a14492 & ~a14474;
assign a14496 = ~a14494 & a14426;
assign a14498 = a14496 & a14420;
assign a14500 = a14498 & a14414;
assign a14502 = a14150 & ~l188;
assign a14504 = a418 & ~i16;
assign a14506 = ~a14504 & ~a14502;
assign a14508 = a14504 & a14502;
assign a14510 = ~a14508 & ~a14506;
assign a14512 = ~a14084 & ~a394;
assign a14514 = a14084 & a394;
assign a14516 = ~a14514 & ~a14512;
assign a14518 = a14516 & a14510;
assign a14520 = a14518 & a14480;
assign a14522 = a14520 & a14486;
assign a14524 = a14522 & a14448;
assign a14526 = a14524 & a14466;
assign a14528 = ~a14152 & ~a420;
assign a14530 = a14152 & a420;
assign a14532 = ~a14530 & ~a14528;
assign a14534 = a14532 & a14516;
assign a14536 = a14534 & a14480;
assign a14538 = a14536 & a14486;
assign a14540 = a14538 & a14448;
assign a14542 = a14540 & a14466;
assign a14544 = ~a14094 & ~a374;
assign a14546 = a14094 & a374;
assign a14548 = ~a14546 & ~a14544;
assign a14550 = a14548 & a14516;
assign a14552 = a14550 & a14480;
assign a14554 = a14552 & a14486;
assign a14556 = a14554 & a14448;
assign a14558 = a14556 & a14466;
assign a14560 = ~a14074 & ~a384;
assign a14562 = a14074 & a384;
assign a14564 = ~a14562 & ~a14560;
assign a14566 = a14564 & a14516;
assign a14568 = a14566 & a14480;
assign a14570 = a14568 & a14486;
assign a14572 = a14570 & a14448;
assign a14574 = a14572 & a14466;
assign a14576 = ~a14102 & ~a402;
assign a14578 = a14102 & a402;
assign a14580 = ~a14578 & ~a14576;
assign a14582 = a14580 & a14516;
assign a14584 = a14582 & a14480;
assign a14586 = a14584 & a14486;
assign a14588 = a14586 & a14448;
assign a14590 = a14588 & a14466;
assign a14592 = ~a14110 & ~a410;
assign a14594 = a14110 & a410;
assign a14596 = ~a14594 & ~a14592;
assign a14598 = a14596 & a14516;
assign a14600 = a14598 & a14480;
assign a14602 = a14600 & a14486;
assign a14604 = a14602 & a14448;
assign a14606 = a14604 & a14466;
assign a14608 = ~a14606 & ~a14590;
assign a14610 = a14608 & ~a14574;
assign a14612 = a14610 & ~a14558;
assign a14614 = a14612 & ~a14542;
assign a14616 = a14614 & ~a14526;
assign a14618 = a14616 & ~a14500;
assign a14620 = ~a14618 & a14408;
assign a14622 = ~l230 & ~i58;
assign a14624 = l230 & i58;
assign a14626 = ~a14624 & ~a14622;
assign a14628 = a14486 & a14430;
assign a14630 = a14628 & a14448;
assign a14632 = a14630 & a14466;
assign a14634 = a14632 & a14426;
assign a14636 = a14634 & a14420;
assign a14638 = a14636 & a14414;
assign a14640 = a14638 & a14626;
assign a14642 = a14632 & a14408;
assign a14644 = a14642 & a14532;
assign a14646 = a14644 & a14510;
assign a14648 = a14548 & a14510;
assign a14650 = a14648 & a14486;
assign a14652 = a14650 & a14430;
assign a14654 = a14652 & a14448;
assign a14656 = a14654 & a14466;
assign a14658 = a14656 & a14408;
assign a14660 = a14548 & a14532;
assign a14662 = a14660 & a14486;
assign a14664 = a14662 & a14430;
assign a14666 = a14664 & a14448;
assign a14668 = a14666 & a14466;
assign a14670 = a14668 & a14408;
assign a14672 = a14564 & a14510;
assign a14674 = a14672 & a14486;
assign a14676 = a14674 & a14430;
assign a14678 = a14676 & a14448;
assign a14680 = a14678 & a14466;
assign a14682 = a14680 & a14408;
assign a14684 = a14564 & a14532;
assign a14686 = a14684 & a14486;
assign a14688 = a14686 & a14430;
assign a14690 = a14688 & a14448;
assign a14692 = a14690 & a14466;
assign a14694 = a14692 & a14408;
assign a14696 = a14564 & a14548;
assign a14698 = a14696 & a14486;
assign a14700 = a14698 & a14430;
assign a14702 = a14700 & a14448;
assign a14704 = a14702 & a14466;
assign a14706 = a14704 & a14408;
assign a14708 = a14580 & a14510;
assign a14710 = a14708 & a14486;
assign a14712 = a14710 & a14430;
assign a14714 = a14712 & a14448;
assign a14716 = a14714 & a14466;
assign a14718 = a14716 & a14408;
assign a14720 = a14580 & a14548;
assign a14722 = a14720 & a14486;
assign a14724 = a14722 & a14430;
assign a14726 = a14724 & a14448;
assign a14728 = a14726 & a14466;
assign a14730 = a14728 & a14408;
assign a14732 = a14580 & a14532;
assign a14734 = a14732 & a14486;
assign a14736 = a14734 & a14430;
assign a14738 = a14736 & a14448;
assign a14740 = a14738 & a14466;
assign a14742 = a14740 & a14408;
assign a14744 = a14580 & a14564;
assign a14746 = a14744 & a14486;
assign a14748 = a14746 & a14430;
assign a14750 = a14748 & a14448;
assign a14752 = a14750 & a14466;
assign a14754 = a14752 & a14408;
assign a14756 = a14596 & a14510;
assign a14758 = a14756 & a14486;
assign a14760 = a14758 & a14430;
assign a14762 = a14760 & a14448;
assign a14764 = a14762 & a14466;
assign a14766 = a14764 & a14408;
assign a14768 = a14596 & a14532;
assign a14770 = a14768 & a14486;
assign a14772 = a14770 & a14430;
assign a14774 = a14772 & a14448;
assign a14776 = a14774 & a14466;
assign a14778 = a14776 & a14408;
assign a14780 = a14596 & a14548;
assign a14782 = a14780 & a14486;
assign a14784 = a14782 & a14430;
assign a14786 = a14784 & a14448;
assign a14788 = a14786 & a14466;
assign a14790 = a14788 & a14408;
assign a14792 = a14596 & a14564;
assign a14794 = a14792 & a14486;
assign a14796 = a14794 & a14430;
assign a14798 = a14796 & a14448;
assign a14800 = a14798 & a14466;
assign a14802 = a14800 & a14408;
assign a14804 = a14596 & a14580;
assign a14806 = a14804 & a14486;
assign a14808 = a14806 & a14430;
assign a14810 = a14808 & a14448;
assign a14812 = a14810 & a14466;
assign a14814 = a14812 & a14408;
assign a14816 = a14642 & a14516;
assign a14818 = a14816 & a14510;
assign a14820 = a14644 & a14516;
assign a14822 = a14642 & a14548;
assign a14824 = a14822 & a14516;
assign a14826 = a14642 & a14564;
assign a14828 = a14826 & a14516;
assign a14830 = a14642 & a14580;
assign a14832 = a14830 & a14516;
assign a14834 = a14642 & a14596;
assign a14836 = a14834 & a14516;
assign a14838 = ~a14836 & ~a14832;
assign a14840 = a14838 & ~a14828;
assign a14842 = a14840 & ~a14824;
assign a14844 = a14842 & ~a14820;
assign a14846 = a14844 & ~a14818;
assign a14848 = a14846 & ~a14814;
assign a14850 = a14848 & ~a14802;
assign a14852 = a14850 & ~a14790;
assign a14854 = a14852 & ~a14778;
assign a14856 = a14854 & ~a14766;
assign a14858 = a14856 & ~a14754;
assign a14860 = a14858 & ~a14742;
assign a14862 = a14860 & ~a14730;
assign a14864 = a14862 & ~a14718;
assign a14866 = a14864 & ~a14706;
assign a14868 = a14866 & ~a14694;
assign a14870 = a14868 & ~a14682;
assign a14872 = a14870 & ~a14670;
assign a14874 = a14872 & ~a14658;
assign a14876 = a14874 & ~a14646;
assign a14878 = a14876 & ~a14640;
assign a14880 = a14878 & ~a14620;
assign a14882 = ~a14880 & a14402;
assign a14884 = ~l226 & ~i54;
assign a14886 = l226 & i54;
assign a14888 = ~a14886 & ~a14884;
assign a14890 = a14642 & a14426;
assign a14892 = a14890 & a14420;
assign a14894 = a14892 & a14414;
assign a14896 = a14894 & a14888;
assign a14898 = ~a14896 & ~a14882;
assign a14900 = ~a14898 & a14396;
assign a14902 = ~l228 & ~i56;
assign a14904 = l228 & i56;
assign a14906 = ~a14904 & ~a14902;
assign a14908 = a14430 & a14402;
assign a14910 = a14908 & a14486;
assign a14912 = a14910 & a14448;
assign a14914 = a14912 & a14466;
assign a14916 = a14914 & a14408;
assign a14918 = a14916 & a14426;
assign a14920 = a14918 & a14420;
assign a14922 = a14920 & a14414;
assign a14924 = a14922 & a14906;
assign a14926 = ~a14924 & ~a14900;
assign a14928 = ~a14926 & a14390;
assign a14930 = ~l224 & ~i52;
assign a14932 = l224 & i52;
assign a14934 = ~a14932 & ~a14930;
assign a14936 = a14430 & a14396;
assign a14938 = a14936 & a14402;
assign a14940 = a14938 & a14486;
assign a14942 = a14940 & a14448;
assign a14944 = a14942 & a14466;
assign a14946 = a14944 & a14408;
assign a14948 = a14946 & a14426;
assign a14950 = a14948 & a14420;
assign a14952 = a14950 & a14414;
assign a14954 = a14952 & a14934;
assign a14956 = ~a14954 & ~a14928;
assign a14958 = ~a14956 & a14384;
assign a14960 = ~l222 & ~i50;
assign a14962 = l222 & i50;
assign a14964 = ~a14962 & ~a14960;
assign a14966 = a14430 & a14390;
assign a14968 = a14966 & a14396;
assign a14970 = a14968 & a14402;
assign a14972 = a14970 & a14486;
assign a14974 = a14972 & a14448;
assign a14976 = a14974 & a14466;
assign a14978 = a14976 & a14408;
assign a14980 = a14978 & a14426;
assign a14982 = a14980 & a14420;
assign a14984 = a14982 & a14414;
assign a14986 = a14984 & a14964;
assign a14988 = ~a14986 & ~a14958;
assign a14990 = ~a14988 & a14378;
assign a14992 = ~l220 & ~i48;
assign a14994 = l220 & i48;
assign a14996 = ~a14994 & ~a14992;
assign a14998 = a14430 & a14384;
assign a15000 = a14998 & a14390;
assign a15002 = a15000 & a14396;
assign a15004 = a15002 & a14402;
assign a15006 = a15004 & a14486;
assign a15008 = a15006 & a14448;
assign a15010 = a15008 & a14466;
assign a15012 = a15010 & a14408;
assign a15014 = a15012 & a14426;
assign a15016 = a15014 & a14420;
assign a15018 = a15016 & a14414;
assign a15020 = a15018 & a14996;
assign a15022 = ~a15020 & ~a14990;
assign a15024 = ~a15022 & a14372;
assign a15026 = a15024 & a14366;
assign a15028 = a15026 & a14360;
assign a15030 = ~a10642 & ~a7938;
assign a15032 = a10642 & a7938;
assign a15034 = ~a15032 & ~a15030;
assign a15036 = ~a7960 & ~a358;
assign a15038 = a7960 & a358;
assign a15040 = ~a15038 & ~a15036;
assign a15042 = a14430 & a14378;
assign a15044 = a15042 & a14384;
assign a15046 = a15044 & a14390;
assign a15048 = a15046 & a14396;
assign a15050 = a15048 & a14402;
assign a15052 = a15050 & a14486;
assign a15054 = a15052 & a14448;
assign a15056 = a15054 & a14466;
assign a15058 = a15056 & a14408;
assign a15060 = a15058 & a14426;
assign a15062 = a15060 & a14420;
assign a15064 = a15062 & a14414;
assign a15066 = a15064 & a15040;
assign a15068 = a15066 & a15034;
assign a15070 = ~a7956 & ~a7950;
assign a15072 = a7956 & a7950;
assign a15074 = ~a15072 & ~a15070;
assign a15076 = a15074 & a15034;
assign a15078 = a15076 & a14378;
assign a15080 = a15078 & a14430;
assign a15082 = a15080 & a14384;
assign a15084 = a15082 & a14390;
assign a15086 = a15084 & a14396;
assign a15088 = a15086 & a14402;
assign a15090 = a15088 & a14486;
assign a15092 = a15090 & a14448;
assign a15094 = a15092 & a14466;
assign a15096 = a15094 & a14408;
assign a15098 = a15096 & a14426;
assign a15100 = a15098 & a14420;
assign a15102 = a15100 & a14414;
assign a15104 = a15074 & a15040;
assign a15106 = a15104 & a14378;
assign a15108 = a15106 & a14430;
assign a15110 = a15108 & a14384;
assign a15112 = a15110 & a14390;
assign a15114 = a15112 & a14396;
assign a15116 = a15114 & a14402;
assign a15118 = a15116 & a14486;
assign a15120 = a15118 & a14448;
assign a15122 = a15120 & a14466;
assign a15124 = a15122 & a14408;
assign a15126 = a15124 & a14426;
assign a15128 = a15126 & a14420;
assign a15130 = a15128 & a14414;
assign a15132 = ~a7932 & ~a354;
assign a15134 = a7932 & a354;
assign a15136 = ~a15134 & ~a15132;
assign a15138 = a15136 & a15034;
assign a15140 = a15138 & a14378;
assign a15142 = a15140 & a14430;
assign a15144 = a15142 & a14384;
assign a15146 = a15144 & a14390;
assign a15148 = a15146 & a14396;
assign a15150 = a15148 & a14402;
assign a15152 = a15150 & a14486;
assign a15154 = a15152 & a14448;
assign a15156 = a15154 & a14466;
assign a15158 = a15156 & a14408;
assign a15160 = a15158 & a14426;
assign a15162 = a15160 & a14420;
assign a15164 = a15162 & a14414;
assign a15166 = a15136 & a15040;
assign a15168 = a15166 & a14378;
assign a15170 = a15168 & a14430;
assign a15172 = a15170 & a14384;
assign a15174 = a15172 & a14390;
assign a15176 = a15174 & a14396;
assign a15178 = a15176 & a14402;
assign a15180 = a15178 & a14486;
assign a15182 = a15180 & a14448;
assign a15184 = a15182 & a14466;
assign a15186 = a15184 & a14408;
assign a15188 = a15186 & a14426;
assign a15190 = a15188 & a14420;
assign a15192 = a15190 & a14414;
assign a15194 = a15136 & a15074;
assign a15196 = a15194 & a14378;
assign a15198 = a15196 & a14430;
assign a15200 = a15198 & a14384;
assign a15202 = a15200 & a14390;
assign a15204 = a15202 & a14396;
assign a15206 = a15204 & a14402;
assign a15208 = a15206 & a14486;
assign a15210 = a15208 & a14448;
assign a15212 = a15210 & a14466;
assign a15214 = a15212 & a14408;
assign a15216 = a15214 & a14426;
assign a15218 = a15216 & a14420;
assign a15220 = a15218 & a14414;
assign a15222 = ~a7928 & ~a7924;
assign a15224 = a7928 & a7924;
assign a15226 = ~a15224 & ~a15222;
assign a15228 = a15226 & a15034;
assign a15230 = a15228 & a14378;
assign a15232 = a15230 & a14430;
assign a15234 = a15232 & a14384;
assign a15236 = a15234 & a14390;
assign a15238 = a15236 & a14396;
assign a15240 = a15238 & a14402;
assign a15242 = a15240 & a14486;
assign a15244 = a15242 & a14448;
assign a15246 = a15244 & a14466;
assign a15248 = a15246 & a14408;
assign a15250 = a15248 & a14426;
assign a15252 = a15250 & a14420;
assign a15254 = a15252 & a14414;
assign a15256 = a15226 & a15040;
assign a15258 = a15256 & a14378;
assign a15260 = a15258 & a14430;
assign a15262 = a15260 & a14384;
assign a15264 = a15262 & a14390;
assign a15266 = a15264 & a14396;
assign a15268 = a15266 & a14402;
assign a15270 = a15268 & a14486;
assign a15272 = a15270 & a14448;
assign a15274 = a15272 & a14466;
assign a15276 = a15274 & a14408;
assign a15278 = a15276 & a14426;
assign a15280 = a15278 & a14420;
assign a15282 = a15280 & a14414;
assign a15284 = a15226 & a15074;
assign a15286 = a15284 & a14378;
assign a15288 = a15286 & a14430;
assign a15290 = a15288 & a14384;
assign a15292 = a15290 & a14390;
assign a15294 = a15292 & a14396;
assign a15296 = a15294 & a14402;
assign a15298 = a15296 & a14486;
assign a15300 = a15298 & a14448;
assign a15302 = a15300 & a14466;
assign a15304 = a15302 & a14408;
assign a15306 = a15304 & a14426;
assign a15308 = a15306 & a14420;
assign a15310 = a15308 & a14414;
assign a15312 = a15226 & a15136;
assign a15314 = a15312 & a14378;
assign a15316 = a15314 & a14430;
assign a15318 = a15316 & a14384;
assign a15320 = a15318 & a14390;
assign a15322 = a15320 & a14396;
assign a15324 = a15322 & a14402;
assign a15326 = a15324 & a14486;
assign a15328 = a15326 & a14448;
assign a15330 = a15328 & a14466;
assign a15332 = a15330 & a14408;
assign a15334 = a15332 & a14426;
assign a15336 = a15334 & a14420;
assign a15338 = a15336 & a14414;
assign a15340 = ~a7606 & ~a6836;
assign a15342 = a7606 & a6836;
assign a15344 = ~a15342 & ~a15340;
assign a15346 = a15344 & a15034;
assign a15348 = a15346 & a14378;
assign a15350 = a15348 & a14430;
assign a15352 = a15350 & a14384;
assign a15354 = a15352 & a14390;
assign a15356 = a15354 & a14396;
assign a15358 = a15356 & a14402;
assign a15360 = a15358 & a14486;
assign a15362 = a15360 & a14448;
assign a15364 = a15362 & a14466;
assign a15366 = a15364 & a14408;
assign a15368 = a15366 & a14426;
assign a15370 = a15368 & a14420;
assign a15372 = a15370 & a14414;
assign a15374 = a15344 & a15040;
assign a15376 = a15374 & a14378;
assign a15378 = a15376 & a14430;
assign a15380 = a15378 & a14384;
assign a15382 = a15380 & a14390;
assign a15384 = a15382 & a14396;
assign a15386 = a15384 & a14402;
assign a15388 = a15386 & a14486;
assign a15390 = a15388 & a14448;
assign a15392 = a15390 & a14466;
assign a15394 = a15392 & a14408;
assign a15396 = a15394 & a14426;
assign a15398 = a15396 & a14420;
assign a15400 = a15398 & a14414;
assign a15402 = a15344 & a15074;
assign a15404 = a15402 & a14378;
assign a15406 = a15404 & a14430;
assign a15408 = a15406 & a14384;
assign a15410 = a15408 & a14390;
assign a15412 = a15410 & a14396;
assign a15414 = a15412 & a14402;
assign a15416 = a15414 & a14486;
assign a15418 = a15416 & a14448;
assign a15420 = a15418 & a14466;
assign a15422 = a15420 & a14408;
assign a15424 = a15422 & a14426;
assign a15426 = a15424 & a14420;
assign a15428 = a15426 & a14414;
assign a15430 = a15344 & a15136;
assign a15432 = a15430 & a14378;
assign a15434 = a15432 & a14430;
assign a15436 = a15434 & a14384;
assign a15438 = a15436 & a14390;
assign a15440 = a15438 & a14396;
assign a15442 = a15440 & a14402;
assign a15444 = a15442 & a14486;
assign a15446 = a15444 & a14448;
assign a15448 = a15446 & a14466;
assign a15450 = a15448 & a14408;
assign a15452 = a15450 & a14426;
assign a15454 = a15452 & a14420;
assign a15456 = a15454 & a14414;
assign a15458 = a15344 & a15226;
assign a15460 = a15458 & a14378;
assign a15462 = a15460 & a14430;
assign a15464 = a15462 & a14384;
assign a15466 = a15464 & a14390;
assign a15468 = a15466 & a14396;
assign a15470 = a15468 & a14402;
assign a15472 = a15470 & a14486;
assign a15474 = a15472 & a14448;
assign a15476 = a15474 & a14466;
assign a15478 = a15476 & a14408;
assign a15480 = a15478 & a14426;
assign a15482 = a15480 & a14420;
assign a15484 = a15482 & a14414;
assign a15486 = a352 & i70;
assign a15488 = ~a15486 & ~a6678;
assign a15490 = a15486 & a6678;
assign a15492 = ~a15490 & ~a15488;
assign a15494 = a15492 & a15034;
assign a15496 = a15494 & a14378;
assign a15498 = a15496 & a14430;
assign a15500 = a15498 & a14384;
assign a15502 = a15500 & a14390;
assign a15504 = a15502 & a14396;
assign a15506 = a15504 & a14402;
assign a15508 = a15506 & a14486;
assign a15510 = a15508 & a14448;
assign a15512 = a15510 & a14466;
assign a15514 = a15512 & a14408;
assign a15516 = a15514 & a14426;
assign a15518 = a15516 & a14420;
assign a15520 = a15518 & a14414;
assign a15522 = a15492 & a15040;
assign a15524 = a15522 & a14378;
assign a15526 = a15524 & a14430;
assign a15528 = a15526 & a14384;
assign a15530 = a15528 & a14390;
assign a15532 = a15530 & a14396;
assign a15534 = a15532 & a14402;
assign a15536 = a15534 & a14486;
assign a15538 = a15536 & a14448;
assign a15540 = a15538 & a14466;
assign a15542 = a15540 & a14408;
assign a15544 = a15542 & a14426;
assign a15546 = a15544 & a14420;
assign a15548 = a15546 & a14414;
assign a15550 = a15492 & a15074;
assign a15552 = a15550 & a14378;
assign a15554 = a15552 & a14430;
assign a15556 = a15554 & a14384;
assign a15558 = a15556 & a14390;
assign a15560 = a15558 & a14396;
assign a15562 = a15560 & a14402;
assign a15564 = a15562 & a14486;
assign a15566 = a15564 & a14448;
assign a15568 = a15566 & a14466;
assign a15570 = a15568 & a14408;
assign a15572 = a15570 & a14426;
assign a15574 = a15572 & a14420;
assign a15576 = a15574 & a14414;
assign a15578 = a15492 & a15136;
assign a15580 = a15578 & a14378;
assign a15582 = a15580 & a14430;
assign a15584 = a15582 & a14384;
assign a15586 = a15584 & a14390;
assign a15588 = a15586 & a14396;
assign a15590 = a15588 & a14402;
assign a15592 = a15590 & a14486;
assign a15594 = a15592 & a14448;
assign a15596 = a15594 & a14466;
assign a15598 = a15596 & a14408;
assign a15600 = a15598 & a14426;
assign a15602 = a15600 & a14420;
assign a15604 = a15602 & a14414;
assign a15606 = a15492 & a15226;
assign a15608 = a15606 & a14378;
assign a15610 = a15608 & a14430;
assign a15612 = a15610 & a14384;
assign a15614 = a15612 & a14390;
assign a15616 = a15614 & a14396;
assign a15618 = a15616 & a14402;
assign a15620 = a15618 & a14486;
assign a15622 = a15620 & a14448;
assign a15624 = a15622 & a14466;
assign a15626 = a15624 & a14408;
assign a15628 = a15626 & a14426;
assign a15630 = a15628 & a14420;
assign a15632 = a15630 & a14414;
assign a15634 = a15492 & a15344;
assign a15636 = a15634 & a14378;
assign a15638 = a15636 & a14430;
assign a15640 = a15638 & a14384;
assign a15642 = a15640 & a14390;
assign a15644 = a15642 & a14396;
assign a15646 = a15644 & a14402;
assign a15648 = a15646 & a14486;
assign a15650 = a15648 & a14448;
assign a15652 = a15650 & a14466;
assign a15654 = a15652 & a14408;
assign a15656 = a15654 & a14426;
assign a15658 = a15656 & a14420;
assign a15660 = a15658 & a14414;
assign a15662 = ~a15660 & ~a15632;
assign a15664 = a15662 & ~a15604;
assign a15666 = a15664 & ~a15576;
assign a15668 = a15666 & ~a15548;
assign a15670 = a15668 & ~a15520;
assign a15672 = a15670 & ~a15484;
assign a15674 = a15672 & ~a15456;
assign a15676 = a15674 & ~a15428;
assign a15678 = a15676 & ~a15400;
assign a15680 = a15678 & ~a15372;
assign a15682 = a15680 & ~a15338;
assign a15684 = a15682 & ~a15310;
assign a15686 = a15684 & ~a15282;
assign a15688 = a15686 & ~a15254;
assign a15690 = a15688 & ~a15220;
assign a15692 = a15690 & ~a15192;
assign a15694 = a15692 & ~a15164;
assign a15696 = a15694 & ~a15130;
assign a15698 = a15696 & ~a15102;
assign a15700 = a15698 & ~a15068;
assign a15702 = a15700 & ~a15028;
assign a15704 = ~a15702 & a14354;
assign a15706 = ~l214 & ~i42;
assign a15708 = l214 & i42;
assign a15710 = ~a15708 & ~a15706;
assign a15712 = a14372 & a14366;
assign a15714 = a15712 & a14360;
assign a15716 = a15714 & a14430;
assign a15718 = a15716 & a14378;
assign a15720 = a15718 & a14384;
assign a15722 = a15720 & a14390;
assign a15724 = a15722 & a14396;
assign a15726 = a15724 & a14402;
assign a15728 = a15726 & a14486;
assign a15730 = a15728 & a14448;
assign a15732 = a15730 & a14466;
assign a15734 = a15732 & a14408;
assign a15736 = a15734 & a14426;
assign a15738 = a15736 & a14420;
assign a15740 = a15738 & a14414;
assign a15742 = a15740 & a15710;
assign a15744 = ~a15742 & ~a15704;
assign a15746 = ~a15744 & a14348;
assign a15748 = ~l212 & ~i40;
assign a15750 = l212 & i40;
assign a15752 = ~a15750 & ~a15748;
assign a15754 = a15716 & a14354;
assign a15756 = a15754 & a14378;
assign a15758 = a15756 & a14384;
assign a15760 = a15758 & a14390;
assign a15762 = a15760 & a14396;
assign a15764 = a15762 & a14402;
assign a15766 = a15764 & a14486;
assign a15768 = a15766 & a14448;
assign a15770 = a15768 & a14466;
assign a15772 = a15770 & a14408;
assign a15774 = a15772 & a14426;
assign a15776 = a15774 & a14420;
assign a15778 = a15776 & a14414;
assign a15780 = a15778 & a15752;
assign a15782 = ~a15780 & ~a15746;
assign a15784 = ~a15782 & a14342;
assign a15786 = ~l210 & ~i38;
assign a15788 = l210 & i38;
assign a15790 = ~a15788 & ~a15786;
assign a15792 = a15716 & a14348;
assign a15794 = a15792 & a14354;
assign a15796 = a15794 & a14378;
assign a15798 = a15796 & a14384;
assign a15800 = a15798 & a14390;
assign a15802 = a15800 & a14396;
assign a15804 = a15802 & a14402;
assign a15806 = a15804 & a14486;
assign a15808 = a15806 & a14448;
assign a15810 = a15808 & a14466;
assign a15812 = a15810 & a14408;
assign a15814 = a15812 & a14426;
assign a15816 = a15814 & a14420;
assign a15818 = a15816 & a14414;
assign a15820 = a15818 & a15790;
assign a15822 = ~a15820 & ~a15784;
assign a15824 = ~a15822 & a14336;
assign a15826 = ~l240 & ~i68;
assign a15828 = l240 & i68;
assign a15830 = ~a15828 & ~a15826;
assign a15832 = a15716 & a14342;
assign a15834 = a15832 & a14348;
assign a15836 = a15834 & a14354;
assign a15838 = a15836 & a14378;
assign a15840 = a15838 & a14384;
assign a15842 = a15840 & a14390;
assign a15844 = a15842 & a14396;
assign a15846 = a15844 & a14402;
assign a15848 = a15846 & a14486;
assign a15850 = a15848 & a14448;
assign a15852 = a15850 & a14466;
assign a15854 = a15852 & a14408;
assign a15856 = a15854 & a14426;
assign a15858 = a15856 & a14420;
assign a15860 = a15858 & a14414;
assign a15862 = a15860 & a15830;
assign a15864 = ~a15862 & ~a15824;
assign a15866 = ~a15864 & a14332;
assign a15868 = ~l208 & ~i36;
assign a15870 = l208 & i36;
assign a15872 = ~a15870 & ~a15868;
assign a15874 = a14430 & a14336;
assign a15876 = a15874 & a14372;
assign a15878 = a15876 & a14366;
assign a15880 = a15878 & a14360;
assign a15882 = a15880 & a14342;
assign a15884 = a15882 & a14348;
assign a15886 = a15884 & a14354;
assign a15888 = a15886 & a14378;
assign a15890 = a15888 & a14384;
assign a15892 = a15890 & a14390;
assign a15894 = a15892 & a14396;
assign a15896 = a15894 & a14402;
assign a15898 = a15896 & a14486;
assign a15900 = a15898 & a14448;
assign a15902 = a15900 & a14466;
assign a15904 = a15902 & a14408;
assign a15906 = a15904 & a14426;
assign a15908 = a15906 & a14420;
assign a15910 = a15908 & a14414;
assign a15912 = a15910 & a15872;
assign a15914 = ~a15912 & ~a15866;
assign a15916 = ~a15914 & a14326;
assign a15918 = ~l232 & ~i60;
assign a15920 = l232 & i60;
assign a15922 = ~a15920 & ~a15918;
assign a15924 = a15880 & a14332;
assign a15926 = a15924 & a14342;
assign a15928 = a15926 & a14348;
assign a15930 = a15928 & a14354;
assign a15932 = a15930 & a14378;
assign a15934 = a15932 & a14384;
assign a15936 = a15934 & a14390;
assign a15938 = a15936 & a14396;
assign a15940 = a15938 & a14402;
assign a15942 = a15940 & a14486;
assign a15944 = a15942 & a14448;
assign a15946 = a15944 & a14466;
assign a15948 = a15946 & a14408;
assign a15950 = a15948 & a14426;
assign a15952 = a15950 & a14420;
assign a15954 = a15952 & a14414;
assign a15956 = a15954 & a15922;
assign a15958 = ~a15956 & ~a15916;
assign a15960 = ~a15958 & a14320;
assign a15962 = ~l264 & ~i92;
assign a15964 = l264 & i92;
assign a15966 = ~a15964 & ~a15962;
assign a15968 = a15880 & a14326;
assign a15970 = a15968 & a14332;
assign a15972 = a15970 & a14342;
assign a15974 = a15972 & a14348;
assign a15976 = a15974 & a14354;
assign a15978 = a15976 & a14378;
assign a15980 = a15978 & a14384;
assign a15982 = a15980 & a14390;
assign a15984 = a15982 & a14396;
assign a15986 = a15984 & a14402;
assign a15988 = a15986 & a14486;
assign a15990 = a15988 & a14448;
assign a15992 = a15990 & a14466;
assign a15994 = a15992 & a14408;
assign a15996 = a15994 & a14426;
assign a15998 = a15996 & a14420;
assign a16000 = a15998 & a14414;
assign a16002 = a16000 & a15966;
assign a16004 = ~a16002 & ~a15960;
assign a16006 = ~a16004 & a14316;
assign a16008 = ~l266 & ~i94;
assign a16010 = l266 & i94;
assign a16012 = ~a16010 & ~a16008;
assign a16014 = a15880 & a14320;
assign a16016 = a16014 & a14326;
assign a16018 = a16016 & a14332;
assign a16020 = a16018 & a14342;
assign a16022 = a16020 & a14348;
assign a16024 = a16022 & a14354;
assign a16026 = a16024 & a14378;
assign a16028 = a16026 & a14384;
assign a16030 = a16028 & a14390;
assign a16032 = a16030 & a14396;
assign a16034 = a16032 & a14402;
assign a16036 = a16034 & a14486;
assign a16038 = a16036 & a14448;
assign a16040 = a16038 & a14466;
assign a16042 = a16040 & a14408;
assign a16044 = a16042 & a14426;
assign a16046 = a16044 & a14420;
assign a16048 = a16046 & a14414;
assign a16050 = a16048 & a16012;
assign a16052 = ~a16050 & ~a16006;
assign a16054 = ~a16052 & a14310;
assign a16056 = a16054 & a14304;
assign a16058 = a16056 & a14298;
assign a16060 = ~a6904 & ~a6898;
assign a16062 = a6904 & a6898;
assign a16064 = ~a16062 & ~a16060;
assign a16066 = ~a7610 & ~a6812;
assign a16068 = a7610 & a6812;
assign a16070 = ~a16068 & ~a16066;
assign a16072 = a15880 & a14316;
assign a16074 = a16072 & a14320;
assign a16076 = a16074 & a14326;
assign a16078 = a16076 & a14332;
assign a16080 = a16078 & a14342;
assign a16082 = a16080 & a14348;
assign a16084 = a16082 & a14354;
assign a16086 = a16084 & a14378;
assign a16088 = a16086 & a14384;
assign a16090 = a16088 & a14390;
assign a16092 = a16090 & a14396;
assign a16094 = a16092 & a14402;
assign a16096 = a16094 & a14486;
assign a16098 = a16096 & a14448;
assign a16100 = a16098 & a14466;
assign a16102 = a16100 & a14408;
assign a16104 = a16102 & a14426;
assign a16106 = a16104 & a14420;
assign a16108 = a16106 & a14414;
assign a16110 = a16108 & a16070;
assign a16112 = a16110 & a16064;
assign a16114 = ~a6884 & ~a6688;
assign a16116 = a6884 & a6688;
assign a16118 = ~a16116 & ~a16114;
assign a16120 = a16118 & a16064;
assign a16122 = a16120 & a14336;
assign a16124 = a16122 & a14430;
assign a16126 = a16124 & a14372;
assign a16128 = a16126 & a14366;
assign a16130 = a16128 & a14360;
assign a16132 = a16130 & a14316;
assign a16134 = a16132 & a14320;
assign a16136 = a16134 & a14326;
assign a16138 = a16136 & a14332;
assign a16140 = a16138 & a14342;
assign a16142 = a16140 & a14348;
assign a16144 = a16142 & a14354;
assign a16146 = a16144 & a14378;
assign a16148 = a16146 & a14384;
assign a16150 = a16148 & a14390;
assign a16152 = a16150 & a14396;
assign a16154 = a16152 & a14402;
assign a16156 = a16154 & a14486;
assign a16158 = a16156 & a14448;
assign a16160 = a16158 & a14466;
assign a16162 = a16160 & a14408;
assign a16164 = a16162 & a14426;
assign a16166 = a16164 & a14420;
assign a16168 = a16166 & a14414;
assign a16170 = a16118 & a16070;
assign a16172 = a16170 & a14336;
assign a16174 = a16172 & a14430;
assign a16176 = a16174 & a14372;
assign a16178 = a16176 & a14366;
assign a16180 = a16178 & a14360;
assign a16182 = a16180 & a14316;
assign a16184 = a16182 & a14320;
assign a16186 = a16184 & a14326;
assign a16188 = a16186 & a14332;
assign a16190 = a16188 & a14342;
assign a16192 = a16190 & a14348;
assign a16194 = a16192 & a14354;
assign a16196 = a16194 & a14378;
assign a16198 = a16196 & a14384;
assign a16200 = a16198 & a14390;
assign a16202 = a16200 & a14396;
assign a16204 = a16202 & a14402;
assign a16206 = a16204 & a14486;
assign a16208 = a16206 & a14448;
assign a16210 = a16208 & a14466;
assign a16212 = a16210 & a14408;
assign a16214 = a16212 & a14426;
assign a16216 = a16214 & a14420;
assign a16218 = a16216 & a14414;
assign a16220 = ~a6976 & ~a6658;
assign a16222 = a6976 & a6658;
assign a16224 = ~a16222 & ~a16220;
assign a16226 = a16224 & a16064;
assign a16228 = a16226 & a14336;
assign a16230 = a16228 & a14430;
assign a16232 = a16230 & a14372;
assign a16234 = a16232 & a14366;
assign a16236 = a16234 & a14360;
assign a16238 = a16236 & a14316;
assign a16240 = a16238 & a14320;
assign a16242 = a16240 & a14326;
assign a16244 = a16242 & a14332;
assign a16246 = a16244 & a14342;
assign a16248 = a16246 & a14348;
assign a16250 = a16248 & a14354;
assign a16252 = a16250 & a14378;
assign a16254 = a16252 & a14384;
assign a16256 = a16254 & a14390;
assign a16258 = a16256 & a14396;
assign a16260 = a16258 & a14402;
assign a16262 = a16260 & a14486;
assign a16264 = a16262 & a14448;
assign a16266 = a16264 & a14466;
assign a16268 = a16266 & a14408;
assign a16270 = a16268 & a14426;
assign a16272 = a16270 & a14420;
assign a16274 = a16272 & a14414;
assign a16276 = a16224 & a16070;
assign a16278 = a16276 & a14336;
assign a16280 = a16278 & a14430;
assign a16282 = a16280 & a14372;
assign a16284 = a16282 & a14366;
assign a16286 = a16284 & a14360;
assign a16288 = a16286 & a14316;
assign a16290 = a16288 & a14320;
assign a16292 = a16290 & a14326;
assign a16294 = a16292 & a14332;
assign a16296 = a16294 & a14342;
assign a16298 = a16296 & a14348;
assign a16300 = a16298 & a14354;
assign a16302 = a16300 & a14378;
assign a16304 = a16302 & a14384;
assign a16306 = a16304 & a14390;
assign a16308 = a16306 & a14396;
assign a16310 = a16308 & a14402;
assign a16312 = a16310 & a14486;
assign a16314 = a16312 & a14448;
assign a16316 = a16314 & a14466;
assign a16318 = a16316 & a14408;
assign a16320 = a16318 & a14426;
assign a16322 = a16320 & a14420;
assign a16324 = a16322 & a14414;
assign a16326 = a16224 & a16118;
assign a16328 = a16326 & a14336;
assign a16330 = a16328 & a14430;
assign a16332 = a16330 & a14372;
assign a16334 = a16332 & a14366;
assign a16336 = a16334 & a14360;
assign a16338 = a16336 & a14316;
assign a16340 = a16338 & a14320;
assign a16342 = a16340 & a14326;
assign a16344 = a16342 & a14332;
assign a16346 = a16344 & a14342;
assign a16348 = a16346 & a14348;
assign a16350 = a16348 & a14354;
assign a16352 = a16350 & a14378;
assign a16354 = a16352 & a14384;
assign a16356 = a16354 & a14390;
assign a16358 = a16356 & a14396;
assign a16360 = a16358 & a14402;
assign a16362 = a16360 & a14486;
assign a16364 = a16362 & a14448;
assign a16366 = a16364 & a14466;
assign a16368 = a16366 & a14408;
assign a16370 = a16368 & a14426;
assign a16372 = a16370 & a14420;
assign a16374 = a16372 & a14414;
assign a16376 = ~a7044 & ~a6730;
assign a16378 = a7044 & a6730;
assign a16380 = ~a16378 & ~a16376;
assign a16382 = a16380 & a16064;
assign a16384 = a16382 & a14336;
assign a16386 = a16384 & a14430;
assign a16388 = a16386 & a14372;
assign a16390 = a16388 & a14366;
assign a16392 = a16390 & a14360;
assign a16394 = a16392 & a14316;
assign a16396 = a16394 & a14320;
assign a16398 = a16396 & a14326;
assign a16400 = a16398 & a14332;
assign a16402 = a16400 & a14342;
assign a16404 = a16402 & a14348;
assign a16406 = a16404 & a14354;
assign a16408 = a16406 & a14378;
assign a16410 = a16408 & a14384;
assign a16412 = a16410 & a14390;
assign a16414 = a16412 & a14396;
assign a16416 = a16414 & a14402;
assign a16418 = a16416 & a14486;
assign a16420 = a16418 & a14448;
assign a16422 = a16420 & a14466;
assign a16424 = a16422 & a14408;
assign a16426 = a16424 & a14426;
assign a16428 = a16426 & a14420;
assign a16430 = a16428 & a14414;
assign a16432 = a16380 & a16070;
assign a16434 = a16432 & a14336;
assign a16436 = a16434 & a14430;
assign a16438 = a16436 & a14372;
assign a16440 = a16438 & a14366;
assign a16442 = a16440 & a14360;
assign a16444 = a16442 & a14316;
assign a16446 = a16444 & a14320;
assign a16448 = a16446 & a14326;
assign a16450 = a16448 & a14332;
assign a16452 = a16450 & a14342;
assign a16454 = a16452 & a14348;
assign a16456 = a16454 & a14354;
assign a16458 = a16456 & a14378;
assign a16460 = a16458 & a14384;
assign a16462 = a16460 & a14390;
assign a16464 = a16462 & a14396;
assign a16466 = a16464 & a14402;
assign a16468 = a16466 & a14486;
assign a16470 = a16468 & a14448;
assign a16472 = a16470 & a14466;
assign a16474 = a16472 & a14408;
assign a16476 = a16474 & a14426;
assign a16478 = a16476 & a14420;
assign a16480 = a16478 & a14414;
assign a16482 = a16380 & a16118;
assign a16484 = a16482 & a14336;
assign a16486 = a16484 & a14430;
assign a16488 = a16486 & a14372;
assign a16490 = a16488 & a14366;
assign a16492 = a16490 & a14360;
assign a16494 = a16492 & a14316;
assign a16496 = a16494 & a14320;
assign a16498 = a16496 & a14326;
assign a16500 = a16498 & a14332;
assign a16502 = a16500 & a14342;
assign a16504 = a16502 & a14348;
assign a16506 = a16504 & a14354;
assign a16508 = a16506 & a14378;
assign a16510 = a16508 & a14384;
assign a16512 = a16510 & a14390;
assign a16514 = a16512 & a14396;
assign a16516 = a16514 & a14402;
assign a16518 = a16516 & a14486;
assign a16520 = a16518 & a14448;
assign a16522 = a16520 & a14466;
assign a16524 = a16522 & a14408;
assign a16526 = a16524 & a14426;
assign a16528 = a16526 & a14420;
assign a16530 = a16528 & a14414;
assign a16532 = a16380 & a16224;
assign a16534 = a16532 & a14336;
assign a16536 = a16534 & a14430;
assign a16538 = a16536 & a14372;
assign a16540 = a16538 & a14366;
assign a16542 = a16540 & a14360;
assign a16544 = a16542 & a14316;
assign a16546 = a16544 & a14320;
assign a16548 = a16546 & a14326;
assign a16550 = a16548 & a14332;
assign a16552 = a16550 & a14342;
assign a16554 = a16552 & a14348;
assign a16556 = a16554 & a14354;
assign a16558 = a16556 & a14378;
assign a16560 = a16558 & a14384;
assign a16562 = a16560 & a14390;
assign a16564 = a16562 & a14396;
assign a16566 = a16564 & a14402;
assign a16568 = a16566 & a14486;
assign a16570 = a16568 & a14448;
assign a16572 = a16570 & a14466;
assign a16574 = a16572 & a14408;
assign a16576 = a16574 & a14426;
assign a16578 = a16576 & a14420;
assign a16580 = a16578 & a14414;
assign a16582 = ~a16580 & ~a16530;
assign a16584 = a16582 & ~a16480;
assign a16586 = a16584 & ~a16430;
assign a16588 = a16586 & ~a16374;
assign a16590 = a16588 & ~a16324;
assign a16592 = a16590 & ~a16274;
assign a16594 = a16592 & ~a16218;
assign a16596 = a16594 & ~a16168;
assign a16598 = a16596 & ~a16112;
assign a16600 = a16598 & ~a16058;
assign a16602 = ~a16600 & a14292;
assign a16604 = ~l262 & ~i90;
assign a16606 = l262 & i90;
assign a16608 = ~a16606 & ~a16604;
assign a16610 = a14310 & a14304;
assign a16612 = a16610 & a14298;
assign a16614 = a16612 & a14430;
assign a16616 = a16614 & a14336;
assign a16618 = a16616 & a14372;
assign a16620 = a16618 & a14366;
assign a16622 = a16620 & a14360;
assign a16624 = a16622 & a14316;
assign a16626 = a16624 & a14320;
assign a16628 = a16626 & a14326;
assign a16630 = a16628 & a14332;
assign a16632 = a16630 & a14342;
assign a16634 = a16632 & a14348;
assign a16636 = a16634 & a14354;
assign a16638 = a16636 & a14378;
assign a16640 = a16638 & a14384;
assign a16642 = a16640 & a14390;
assign a16644 = a16642 & a14396;
assign a16646 = a16644 & a14402;
assign a16648 = a16646 & a14486;
assign a16650 = a16648 & a14448;
assign a16652 = a16650 & a14466;
assign a16654 = a16652 & a14408;
assign a16656 = a16654 & a14426;
assign a16658 = a16656 & a14420;
assign a16660 = a16658 & a14414;
assign a16662 = a16660 & a16608;
assign a16664 = ~a16662 & ~a16602;
assign a16666 = ~a16664 & a14288;
assign a16668 = ~l260 & ~i88;
assign a16670 = l260 & i88;
assign a16672 = ~a16670 & ~a16668;
assign a16674 = a14430 & a14292;
assign a16676 = a16674 & a14310;
assign a16678 = a16676 & a14304;
assign a16680 = a16678 & a14298;
assign a16682 = a16680 & a14336;
assign a16684 = a16682 & a14372;
assign a16686 = a16684 & a14366;
assign a16688 = a16686 & a14360;
assign a16690 = a16688 & a14316;
assign a16692 = a16690 & a14320;
assign a16694 = a16692 & a14326;
assign a16696 = a16694 & a14332;
assign a16698 = a16696 & a14342;
assign a16700 = a16698 & a14348;
assign a16702 = a16700 & a14354;
assign a16704 = a16702 & a14378;
assign a16706 = a16704 & a14384;
assign a16708 = a16706 & a14390;
assign a16710 = a16708 & a14396;
assign a16712 = a16710 & a14402;
assign a16714 = a16712 & a14486;
assign a16716 = a16714 & a14448;
assign a16718 = a16716 & a14466;
assign a16720 = a16718 & a14408;
assign a16722 = a16720 & a14426;
assign a16724 = a16722 & a14420;
assign a16726 = a16724 & a14414;
assign a16728 = a16726 & a16672;
assign a16730 = ~a16728 & ~a16666;
assign a16732 = ~a16730 & a14284;
assign a16734 = ~l308 & ~i136;
assign a16736 = l308 & i136;
assign a16738 = ~a16736 & ~a16734;
assign a16740 = a14430 & a14288;
assign a16742 = a16740 & a14292;
assign a16744 = a16742 & a14310;
assign a16746 = a16744 & a14304;
assign a16748 = a16746 & a14298;
assign a16750 = a16748 & a14336;
assign a16752 = a16750 & a14372;
assign a16754 = a16752 & a14366;
assign a16756 = a16754 & a14360;
assign a16758 = a16756 & a14316;
assign a16760 = a16758 & a14320;
assign a16762 = a16760 & a14326;
assign a16764 = a16762 & a14332;
assign a16766 = a16764 & a14342;
assign a16768 = a16766 & a14348;
assign a16770 = a16768 & a14354;
assign a16772 = a16770 & a14378;
assign a16774 = a16772 & a14384;
assign a16776 = a16774 & a14390;
assign a16778 = a16776 & a14396;
assign a16780 = a16778 & a14402;
assign a16782 = a16780 & a14486;
assign a16784 = a16782 & a14448;
assign a16786 = a16784 & a14466;
assign a16788 = a16786 & a14408;
assign a16790 = a16788 & a14426;
assign a16792 = a16790 & a14420;
assign a16794 = a16792 & a14414;
assign a16796 = a16794 & a16738;
assign a16798 = ~a16796 & ~a16732;
assign a16800 = ~a16798 & a14278;
assign a16802 = ~l306 & ~i134;
assign a16804 = l306 & i134;
assign a16806 = ~a16804 & ~a16802;
assign a16808 = a14430 & a14284;
assign a16810 = a16808 & a14288;
assign a16812 = a16810 & a14292;
assign a16814 = a16812 & a14310;
assign a16816 = a16814 & a14304;
assign a16818 = a16816 & a14298;
assign a16820 = a16818 & a14336;
assign a16822 = a16820 & a14372;
assign a16824 = a16822 & a14366;
assign a16826 = a16824 & a14360;
assign a16828 = a16826 & a14316;
assign a16830 = a16828 & a14320;
assign a16832 = a16830 & a14326;
assign a16834 = a16832 & a14332;
assign a16836 = a16834 & a14342;
assign a16838 = a16836 & a14348;
assign a16840 = a16838 & a14354;
assign a16842 = a16840 & a14378;
assign a16844 = a16842 & a14384;
assign a16846 = a16844 & a14390;
assign a16848 = a16846 & a14396;
assign a16850 = a16848 & a14402;
assign a16852 = a16850 & a14486;
assign a16854 = a16852 & a14448;
assign a16856 = a16854 & a14466;
assign a16858 = a16856 & a14408;
assign a16860 = a16858 & a14426;
assign a16862 = a16860 & a14420;
assign a16864 = a16862 & a14414;
assign a16866 = a16864 & a16806;
assign a16868 = ~a16866 & ~a16800;
assign a16870 = ~a16868 & a14272;
assign a16872 = ~l304 & ~i132;
assign a16874 = l304 & i132;
assign a16876 = ~a16874 & ~a16872;
assign a16878 = a14284 & a14278;
assign a16880 = a16878 & a14430;
assign a16882 = a16880 & a14288;
assign a16884 = a16882 & a14292;
assign a16886 = a16884 & a14310;
assign a16888 = a16886 & a14304;
assign a16890 = a16888 & a14298;
assign a16892 = a16890 & a14336;
assign a16894 = a16892 & a14372;
assign a16896 = a16894 & a14366;
assign a16898 = a16896 & a14360;
assign a16900 = a16898 & a14316;
assign a16902 = a16900 & a14320;
assign a16904 = a16902 & a14326;
assign a16906 = a16904 & a14332;
assign a16908 = a16906 & a14342;
assign a16910 = a16908 & a14348;
assign a16912 = a16910 & a14354;
assign a16914 = a16912 & a14378;
assign a16916 = a16914 & a14384;
assign a16918 = a16916 & a14390;
assign a16920 = a16918 & a14396;
assign a16922 = a16920 & a14402;
assign a16924 = a16922 & a14486;
assign a16926 = a16924 & a14448;
assign a16928 = a16926 & a14466;
assign a16930 = a16928 & a14408;
assign a16932 = a16930 & a14426;
assign a16934 = a16932 & a14420;
assign a16936 = a16934 & a14414;
assign a16938 = a16936 & a16876;
assign a16940 = ~a16938 & ~a16870;
assign a16942 = ~a16940 & a14266;
assign a16944 = ~l302 & ~i130;
assign a16946 = l302 & i130;
assign a16948 = ~a16946 & ~a16944;
assign a16950 = a14278 & a14272;
assign a16952 = a16950 & a14284;
assign a16954 = a16952 & a14430;
assign a16956 = a16954 & a14288;
assign a16958 = a16956 & a14292;
assign a16960 = a16958 & a14310;
assign a16962 = a16960 & a14304;
assign a16964 = a16962 & a14298;
assign a16966 = a16964 & a14336;
assign a16968 = a16966 & a14372;
assign a16970 = a16968 & a14366;
assign a16972 = a16970 & a14360;
assign a16974 = a16972 & a14316;
assign a16976 = a16974 & a14320;
assign a16978 = a16976 & a14326;
assign a16980 = a16978 & a14332;
assign a16982 = a16980 & a14342;
assign a16984 = a16982 & a14348;
assign a16986 = a16984 & a14354;
assign a16988 = a16986 & a14378;
assign a16990 = a16988 & a14384;
assign a16992 = a16990 & a14390;
assign a16994 = a16992 & a14396;
assign a16996 = a16994 & a14402;
assign a16998 = a16996 & a14486;
assign a17000 = a16998 & a14448;
assign a17002 = a17000 & a14466;
assign a17004 = a17002 & a14408;
assign a17006 = a17004 & a14426;
assign a17008 = a17006 & a14420;
assign a17010 = a17008 & a14414;
assign a17012 = a17010 & a16948;
assign a17014 = ~a17012 & ~a16942;
assign a17016 = ~a17014 & a14260;
assign a17018 = ~l292 & ~i120;
assign a17020 = l292 & i120;
assign a17022 = ~a17020 & ~a17018;
assign a17024 = a14272 & a14266;
assign a17026 = a17024 & a14278;
assign a17028 = a17026 & a14284;
assign a17030 = a17028 & a14430;
assign a17032 = a17030 & a14288;
assign a17034 = a17032 & a14292;
assign a17036 = a17034 & a14310;
assign a17038 = a17036 & a14304;
assign a17040 = a17038 & a14298;
assign a17042 = a17040 & a14336;
assign a17044 = a17042 & a14372;
assign a17046 = a17044 & a14366;
assign a17048 = a17046 & a14360;
assign a17050 = a17048 & a14316;
assign a17052 = a17050 & a14320;
assign a17054 = a17052 & a14326;
assign a17056 = a17054 & a14332;
assign a17058 = a17056 & a14342;
assign a17060 = a17058 & a14348;
assign a17062 = a17060 & a14354;
assign a17064 = a17062 & a14378;
assign a17066 = a17064 & a14384;
assign a17068 = a17066 & a14390;
assign a17070 = a17068 & a14396;
assign a17072 = a17070 & a14402;
assign a17074 = a17072 & a14486;
assign a17076 = a17074 & a14448;
assign a17078 = a17076 & a14466;
assign a17080 = a17078 & a14408;
assign a17082 = a17080 & a14426;
assign a17084 = a17082 & a14420;
assign a17086 = a17084 & a14414;
assign a17088 = a17086 & a17022;
assign a17090 = ~a17088 & ~a17016;
assign a17092 = ~a17090 & a14254;
assign a17094 = ~l294 & ~i122;
assign a17096 = l294 & i122;
assign a17098 = ~a17096 & ~a17094;
assign a17100 = a14266 & a14260;
assign a17102 = a17100 & a14272;
assign a17104 = a17102 & a14278;
assign a17106 = a17104 & a14284;
assign a17108 = a17106 & a14430;
assign a17110 = a17108 & a14288;
assign a17112 = a17110 & a14292;
assign a17114 = a17112 & a14310;
assign a17116 = a17114 & a14304;
assign a17118 = a17116 & a14298;
assign a17120 = a17118 & a14336;
assign a17122 = a17120 & a14372;
assign a17124 = a17122 & a14366;
assign a17126 = a17124 & a14360;
assign a17128 = a17126 & a14316;
assign a17130 = a17128 & a14320;
assign a17132 = a17130 & a14326;
assign a17134 = a17132 & a14332;
assign a17136 = a17134 & a14342;
assign a17138 = a17136 & a14348;
assign a17140 = a17138 & a14354;
assign a17142 = a17140 & a14378;
assign a17144 = a17142 & a14384;
assign a17146 = a17144 & a14390;
assign a17148 = a17146 & a14396;
assign a17150 = a17148 & a14402;
assign a17152 = a17150 & a14486;
assign a17154 = a17152 & a14448;
assign a17156 = a17154 & a14466;
assign a17158 = a17156 & a14408;
assign a17160 = a17158 & a14426;
assign a17162 = a17160 & a14420;
assign a17164 = a17162 & a14414;
assign a17166 = a17164 & a17098;
assign a17168 = ~a17166 & ~a17092;
assign a17170 = ~a17168 & a14248;
assign a17172 = ~l300 & ~i128;
assign a17174 = l300 & i128;
assign a17176 = ~a17174 & ~a17172;
assign a17178 = a14260 & a14254;
assign a17180 = a17178 & a14266;
assign a17182 = a17180 & a14272;
assign a17184 = a17182 & a14278;
assign a17186 = a17184 & a14284;
assign a17188 = a17186 & a14430;
assign a17190 = a17188 & a14288;
assign a17192 = a17190 & a14292;
assign a17194 = a17192 & a14310;
assign a17196 = a17194 & a14304;
assign a17198 = a17196 & a14298;
assign a17200 = a17198 & a14336;
assign a17202 = a17200 & a14372;
assign a17204 = a17202 & a14366;
assign a17206 = a17204 & a14360;
assign a17208 = a17206 & a14316;
assign a17210 = a17208 & a14320;
assign a17212 = a17210 & a14326;
assign a17214 = a17212 & a14332;
assign a17216 = a17214 & a14342;
assign a17218 = a17216 & a14348;
assign a17220 = a17218 & a14354;
assign a17222 = a17220 & a14378;
assign a17224 = a17222 & a14384;
assign a17226 = a17224 & a14390;
assign a17228 = a17226 & a14396;
assign a17230 = a17228 & a14402;
assign a17232 = a17230 & a14486;
assign a17234 = a17232 & a14448;
assign a17236 = a17234 & a14466;
assign a17238 = a17236 & a14408;
assign a17240 = a17238 & a14426;
assign a17242 = a17240 & a14420;
assign a17244 = a17242 & a14414;
assign a17246 = a17244 & a17176;
assign a17248 = ~a17246 & ~a17170;
assign a17250 = ~a17248 & a14242;
assign a17252 = ~l298 & ~i126;
assign a17254 = l298 & i126;
assign a17256 = ~a17254 & ~a17252;
assign a17258 = a14254 & a14248;
assign a17260 = a17258 & a14260;
assign a17262 = a17260 & a14266;
assign a17264 = a17262 & a14272;
assign a17266 = a17264 & a14278;
assign a17268 = a17266 & a14284;
assign a17270 = a17268 & a14430;
assign a17272 = a17270 & a14288;
assign a17274 = a17272 & a14292;
assign a17276 = a17274 & a14310;
assign a17278 = a17276 & a14304;
assign a17280 = a17278 & a14298;
assign a17282 = a17280 & a14336;
assign a17284 = a17282 & a14372;
assign a17286 = a17284 & a14366;
assign a17288 = a17286 & a14360;
assign a17290 = a17288 & a14316;
assign a17292 = a17290 & a14320;
assign a17294 = a17292 & a14326;
assign a17296 = a17294 & a14332;
assign a17298 = a17296 & a14342;
assign a17300 = a17298 & a14348;
assign a17302 = a17300 & a14354;
assign a17304 = a17302 & a14378;
assign a17306 = a17304 & a14384;
assign a17308 = a17306 & a14390;
assign a17310 = a17308 & a14396;
assign a17312 = a17310 & a14402;
assign a17314 = a17312 & a14486;
assign a17316 = a17314 & a14448;
assign a17318 = a17316 & a14466;
assign a17320 = a17318 & a14408;
assign a17322 = a17320 & a14426;
assign a17324 = a17322 & a14420;
assign a17326 = a17324 & a14414;
assign a17328 = a17326 & a17256;
assign a17330 = ~a17328 & ~a17250;
assign a17332 = ~a17330 & a14238;
assign a17334 = ~l296 & ~i124;
assign a17336 = l296 & i124;
assign a17338 = ~a17336 & ~a17334;
assign a17340 = a17326 & a14242;
assign a17342 = a17340 & a17338;
assign a17344 = ~a17342 & ~a17332;
assign a17346 = ~a17344 & a14232;
assign a17348 = a17346 & a14226;
assign a17350 = a17348 & a14220;
assign a17352 = a1082 & l278;
assign a17354 = a430 & i106;
assign a17356 = ~a17354 & ~a17352;
assign a17358 = a17354 & a17352;
assign a17360 = ~a17358 & ~a17356;
assign a17362 = ~a952 & ~a438;
assign a17364 = a952 & a438;
assign a17366 = ~a17364 & ~a17362;
assign a17368 = a14254 & a14238;
assign a17370 = a17368 & a14248;
assign a17372 = a17370 & a14260;
assign a17374 = a17372 & a14266;
assign a17376 = a17374 & a14272;
assign a17378 = a17376 & a14278;
assign a17380 = a17378 & a14284;
assign a17382 = a17380 & a14430;
assign a17384 = a17382 & a14288;
assign a17386 = a17384 & a14292;
assign a17388 = a17386 & a14310;
assign a17390 = a17388 & a14304;
assign a17392 = a17390 & a14298;
assign a17394 = a17392 & a14336;
assign a17396 = a17394 & a14372;
assign a17398 = a17396 & a14366;
assign a17400 = a17398 & a14360;
assign a17402 = a17400 & a14316;
assign a17404 = a17402 & a14320;
assign a17406 = a17404 & a14326;
assign a17408 = a17406 & a14332;
assign a17410 = a17408 & a14342;
assign a17412 = a17410 & a14348;
assign a17414 = a17412 & a14354;
assign a17416 = a17414 & a14378;
assign a17418 = a17416 & a14384;
assign a17420 = a17418 & a14390;
assign a17422 = a17420 & a14396;
assign a17424 = a17422 & a14402;
assign a17426 = a17424 & a14486;
assign a17428 = a17426 & a14448;
assign a17430 = a17428 & a14466;
assign a17432 = a17430 & a14408;
assign a17434 = a17432 & a14426;
assign a17436 = a17434 & a14420;
assign a17438 = a17436 & a14414;
assign a17440 = a17438 & a14242;
assign a17442 = a17440 & a17366;
assign a17444 = a17442 & a17360;
assign a17446 = ~a960 & ~a466;
assign a17448 = a960 & a466;
assign a17450 = ~a17448 & ~a17446;
assign a17452 = a17450 & a17360;
assign a17454 = a17452 & a14238;
assign a17456 = a17454 & a14254;
assign a17458 = a17456 & a14248;
assign a17460 = a17458 & a14260;
assign a17462 = a17460 & a14266;
assign a17464 = a17462 & a14272;
assign a17466 = a17464 & a14278;
assign a17468 = a17466 & a14284;
assign a17470 = a17468 & a14430;
assign a17472 = a17470 & a14288;
assign a17474 = a17472 & a14292;
assign a17476 = a17474 & a14310;
assign a17478 = a17476 & a14304;
assign a17480 = a17478 & a14298;
assign a17482 = a17480 & a14336;
assign a17484 = a17482 & a14372;
assign a17486 = a17484 & a14366;
assign a17488 = a17486 & a14360;
assign a17490 = a17488 & a14316;
assign a17492 = a17490 & a14320;
assign a17494 = a17492 & a14326;
assign a17496 = a17494 & a14332;
assign a17498 = a17496 & a14342;
assign a17500 = a17498 & a14348;
assign a17502 = a17500 & a14354;
assign a17504 = a17502 & a14378;
assign a17506 = a17504 & a14384;
assign a17508 = a17506 & a14390;
assign a17510 = a17508 & a14396;
assign a17512 = a17510 & a14402;
assign a17514 = a17512 & a14486;
assign a17516 = a17514 & a14448;
assign a17518 = a17516 & a14466;
assign a17520 = a17518 & a14408;
assign a17522 = a17520 & a14426;
assign a17524 = a17522 & a14420;
assign a17526 = a17524 & a14414;
assign a17528 = a17526 & a14242;
assign a17530 = a17450 & a17366;
assign a17532 = a17530 & a14238;
assign a17534 = a17532 & a14254;
assign a17536 = a17534 & a14248;
assign a17538 = a17536 & a14260;
assign a17540 = a17538 & a14266;
assign a17542 = a17540 & a14272;
assign a17544 = a17542 & a14278;
assign a17546 = a17544 & a14284;
assign a17548 = a17546 & a14430;
assign a17550 = a17548 & a14288;
assign a17552 = a17550 & a14292;
assign a17554 = a17552 & a14310;
assign a17556 = a17554 & a14304;
assign a17558 = a17556 & a14298;
assign a17560 = a17558 & a14336;
assign a17562 = a17560 & a14372;
assign a17564 = a17562 & a14366;
assign a17566 = a17564 & a14360;
assign a17568 = a17566 & a14316;
assign a17570 = a17568 & a14320;
assign a17572 = a17570 & a14326;
assign a17574 = a17572 & a14332;
assign a17576 = a17574 & a14342;
assign a17578 = a17576 & a14348;
assign a17580 = a17578 & a14354;
assign a17582 = a17580 & a14378;
assign a17584 = a17582 & a14384;
assign a17586 = a17584 & a14390;
assign a17588 = a17586 & a14396;
assign a17590 = a17588 & a14402;
assign a17592 = a17590 & a14486;
assign a17594 = a17592 & a14448;
assign a17596 = a17594 & a14466;
assign a17598 = a17596 & a14408;
assign a17600 = a17598 & a14426;
assign a17602 = a17600 & a14420;
assign a17604 = a17602 & a14414;
assign a17606 = a17604 & a14242;
assign a17608 = ~a864 & ~a444;
assign a17610 = a864 & a444;
assign a17612 = ~a17610 & ~a17608;
assign a17614 = a17612 & a17360;
assign a17616 = a17614 & a14238;
assign a17618 = a17616 & a14254;
assign a17620 = a17618 & a14248;
assign a17622 = a17620 & a14260;
assign a17624 = a17622 & a14266;
assign a17626 = a17624 & a14272;
assign a17628 = a17626 & a14278;
assign a17630 = a17628 & a14284;
assign a17632 = a17630 & a14430;
assign a17634 = a17632 & a14288;
assign a17636 = a17634 & a14292;
assign a17638 = a17636 & a14310;
assign a17640 = a17638 & a14304;
assign a17642 = a17640 & a14298;
assign a17644 = a17642 & a14336;
assign a17646 = a17644 & a14372;
assign a17648 = a17646 & a14366;
assign a17650 = a17648 & a14360;
assign a17652 = a17650 & a14316;
assign a17654 = a17652 & a14320;
assign a17656 = a17654 & a14326;
assign a17658 = a17656 & a14332;
assign a17660 = a17658 & a14342;
assign a17662 = a17660 & a14348;
assign a17664 = a17662 & a14354;
assign a17666 = a17664 & a14378;
assign a17668 = a17666 & a14384;
assign a17670 = a17668 & a14390;
assign a17672 = a17670 & a14396;
assign a17674 = a17672 & a14402;
assign a17676 = a17674 & a14486;
assign a17678 = a17676 & a14448;
assign a17680 = a17678 & a14466;
assign a17682 = a17680 & a14408;
assign a17684 = a17682 & a14426;
assign a17686 = a17684 & a14420;
assign a17688 = a17686 & a14414;
assign a17690 = a17688 & a14242;
assign a17692 = a17612 & a17366;
assign a17694 = a17692 & a14238;
assign a17696 = a17694 & a14254;
assign a17698 = a17696 & a14248;
assign a17700 = a17698 & a14260;
assign a17702 = a17700 & a14266;
assign a17704 = a17702 & a14272;
assign a17706 = a17704 & a14278;
assign a17708 = a17706 & a14284;
assign a17710 = a17708 & a14430;
assign a17712 = a17710 & a14288;
assign a17714 = a17712 & a14292;
assign a17716 = a17714 & a14310;
assign a17718 = a17716 & a14304;
assign a17720 = a17718 & a14298;
assign a17722 = a17720 & a14336;
assign a17724 = a17722 & a14372;
assign a17726 = a17724 & a14366;
assign a17728 = a17726 & a14360;
assign a17730 = a17728 & a14316;
assign a17732 = a17730 & a14320;
assign a17734 = a17732 & a14326;
assign a17736 = a17734 & a14332;
assign a17738 = a17736 & a14342;
assign a17740 = a17738 & a14348;
assign a17742 = a17740 & a14354;
assign a17744 = a17742 & a14378;
assign a17746 = a17744 & a14384;
assign a17748 = a17746 & a14390;
assign a17750 = a17748 & a14396;
assign a17752 = a17750 & a14402;
assign a17754 = a17752 & a14486;
assign a17756 = a17754 & a14448;
assign a17758 = a17756 & a14466;
assign a17760 = a17758 & a14408;
assign a17762 = a17760 & a14426;
assign a17764 = a17762 & a14420;
assign a17766 = a17764 & a14414;
assign a17768 = a17766 & a14242;
assign a17770 = a17612 & a17450;
assign a17772 = a17770 & a14238;
assign a17774 = a17772 & a14254;
assign a17776 = a17774 & a14248;
assign a17778 = a17776 & a14260;
assign a17780 = a17778 & a14266;
assign a17782 = a17780 & a14272;
assign a17784 = a17782 & a14278;
assign a17786 = a17784 & a14284;
assign a17788 = a17786 & a14430;
assign a17790 = a17788 & a14288;
assign a17792 = a17790 & a14292;
assign a17794 = a17792 & a14310;
assign a17796 = a17794 & a14304;
assign a17798 = a17796 & a14298;
assign a17800 = a17798 & a14336;
assign a17802 = a17800 & a14372;
assign a17804 = a17802 & a14366;
assign a17806 = a17804 & a14360;
assign a17808 = a17806 & a14316;
assign a17810 = a17808 & a14320;
assign a17812 = a17810 & a14326;
assign a17814 = a17812 & a14332;
assign a17816 = a17814 & a14342;
assign a17818 = a17816 & a14348;
assign a17820 = a17818 & a14354;
assign a17822 = a17820 & a14378;
assign a17824 = a17822 & a14384;
assign a17826 = a17824 & a14390;
assign a17828 = a17826 & a14396;
assign a17830 = a17828 & a14402;
assign a17832 = a17830 & a14486;
assign a17834 = a17832 & a14448;
assign a17836 = a17834 & a14466;
assign a17838 = a17836 & a14408;
assign a17840 = a17838 & a14426;
assign a17842 = a17840 & a14420;
assign a17844 = a17842 & a14414;
assign a17846 = a17844 & a14242;
assign a17848 = ~a1062 & ~a448;
assign a17850 = a1062 & a448;
assign a17852 = ~a17850 & ~a17848;
assign a17854 = a17852 & a17360;
assign a17856 = a17854 & a14238;
assign a17858 = a17856 & a14254;
assign a17860 = a17858 & a14248;
assign a17862 = a17860 & a14260;
assign a17864 = a17862 & a14266;
assign a17866 = a17864 & a14272;
assign a17868 = a17866 & a14278;
assign a17870 = a17868 & a14284;
assign a17872 = a17870 & a14430;
assign a17874 = a17872 & a14288;
assign a17876 = a17874 & a14292;
assign a17878 = a17876 & a14310;
assign a17880 = a17878 & a14304;
assign a17882 = a17880 & a14298;
assign a17884 = a17882 & a14336;
assign a17886 = a17884 & a14372;
assign a17888 = a17886 & a14366;
assign a17890 = a17888 & a14360;
assign a17892 = a17890 & a14316;
assign a17894 = a17892 & a14320;
assign a17896 = a17894 & a14326;
assign a17898 = a17896 & a14332;
assign a17900 = a17898 & a14342;
assign a17902 = a17900 & a14348;
assign a17904 = a17902 & a14354;
assign a17906 = a17904 & a14378;
assign a17908 = a17906 & a14384;
assign a17910 = a17908 & a14390;
assign a17912 = a17910 & a14396;
assign a17914 = a17912 & a14402;
assign a17916 = a17914 & a14486;
assign a17918 = a17916 & a14448;
assign a17920 = a17918 & a14466;
assign a17922 = a17920 & a14408;
assign a17924 = a17922 & a14426;
assign a17926 = a17924 & a14420;
assign a17928 = a17926 & a14414;
assign a17930 = a17928 & a14242;
assign a17932 = a17852 & a17366;
assign a17934 = a17932 & a14238;
assign a17936 = a17934 & a14254;
assign a17938 = a17936 & a14248;
assign a17940 = a17938 & a14260;
assign a17942 = a17940 & a14266;
assign a17944 = a17942 & a14272;
assign a17946 = a17944 & a14278;
assign a17948 = a17946 & a14284;
assign a17950 = a17948 & a14430;
assign a17952 = a17950 & a14288;
assign a17954 = a17952 & a14292;
assign a17956 = a17954 & a14310;
assign a17958 = a17956 & a14304;
assign a17960 = a17958 & a14298;
assign a17962 = a17960 & a14336;
assign a17964 = a17962 & a14372;
assign a17966 = a17964 & a14366;
assign a17968 = a17966 & a14360;
assign a17970 = a17968 & a14316;
assign a17972 = a17970 & a14320;
assign a17974 = a17972 & a14326;
assign a17976 = a17974 & a14332;
assign a17978 = a17976 & a14342;
assign a17980 = a17978 & a14348;
assign a17982 = a17980 & a14354;
assign a17984 = a17982 & a14378;
assign a17986 = a17984 & a14384;
assign a17988 = a17986 & a14390;
assign a17990 = a17988 & a14396;
assign a17992 = a17990 & a14402;
assign a17994 = a17992 & a14486;
assign a17996 = a17994 & a14448;
assign a17998 = a17996 & a14466;
assign a18000 = a17998 & a14408;
assign a18002 = a18000 & a14426;
assign a18004 = a18002 & a14420;
assign a18006 = a18004 & a14414;
assign a18008 = a18006 & a14242;
assign a18010 = a17852 & a17450;
assign a18012 = a18010 & a14238;
assign a18014 = a18012 & a14254;
assign a18016 = a18014 & a14248;
assign a18018 = a18016 & a14260;
assign a18020 = a18018 & a14266;
assign a18022 = a18020 & a14272;
assign a18024 = a18022 & a14278;
assign a18026 = a18024 & a14284;
assign a18028 = a18026 & a14430;
assign a18030 = a18028 & a14288;
assign a18032 = a18030 & a14292;
assign a18034 = a18032 & a14310;
assign a18036 = a18034 & a14304;
assign a18038 = a18036 & a14298;
assign a18040 = a18038 & a14336;
assign a18042 = a18040 & a14372;
assign a18044 = a18042 & a14366;
assign a18046 = a18044 & a14360;
assign a18048 = a18046 & a14316;
assign a18050 = a18048 & a14320;
assign a18052 = a18050 & a14326;
assign a18054 = a18052 & a14332;
assign a18056 = a18054 & a14342;
assign a18058 = a18056 & a14348;
assign a18060 = a18058 & a14354;
assign a18062 = a18060 & a14378;
assign a18064 = a18062 & a14384;
assign a18066 = a18064 & a14390;
assign a18068 = a18066 & a14396;
assign a18070 = a18068 & a14402;
assign a18072 = a18070 & a14486;
assign a18074 = a18072 & a14448;
assign a18076 = a18074 & a14466;
assign a18078 = a18076 & a14408;
assign a18080 = a18078 & a14426;
assign a18082 = a18080 & a14420;
assign a18084 = a18082 & a14414;
assign a18086 = a18084 & a14242;
assign a18088 = a17852 & a17612;
assign a18090 = a18088 & a14238;
assign a18092 = a18090 & a14254;
assign a18094 = a18092 & a14248;
assign a18096 = a18094 & a14260;
assign a18098 = a18096 & a14266;
assign a18100 = a18098 & a14272;
assign a18102 = a18100 & a14278;
assign a18104 = a18102 & a14284;
assign a18106 = a18104 & a14430;
assign a18108 = a18106 & a14288;
assign a18110 = a18108 & a14292;
assign a18112 = a18110 & a14310;
assign a18114 = a18112 & a14304;
assign a18116 = a18114 & a14298;
assign a18118 = a18116 & a14336;
assign a18120 = a18118 & a14372;
assign a18122 = a18120 & a14366;
assign a18124 = a18122 & a14360;
assign a18126 = a18124 & a14316;
assign a18128 = a18126 & a14320;
assign a18130 = a18128 & a14326;
assign a18132 = a18130 & a14332;
assign a18134 = a18132 & a14342;
assign a18136 = a18134 & a14348;
assign a18138 = a18136 & a14354;
assign a18140 = a18138 & a14378;
assign a18142 = a18140 & a14384;
assign a18144 = a18142 & a14390;
assign a18146 = a18144 & a14396;
assign a18148 = a18146 & a14402;
assign a18150 = a18148 & a14486;
assign a18152 = a18150 & a14448;
assign a18154 = a18152 & a14466;
assign a18156 = a18154 & a14408;
assign a18158 = a18156 & a14426;
assign a18160 = a18158 & a14420;
assign a18162 = a18160 & a14414;
assign a18164 = a18162 & a14242;
assign a18166 = ~a1084 & ~a432;
assign a18168 = a1084 & a432;
assign a18170 = ~a18168 & ~a18166;
assign a18172 = a18170 & a17360;
assign a18174 = a18172 & a14238;
assign a18176 = a18174 & a14254;
assign a18178 = a18176 & a14248;
assign a18180 = a18178 & a14260;
assign a18182 = a18180 & a14266;
assign a18184 = a18182 & a14272;
assign a18186 = a18184 & a14278;
assign a18188 = a18186 & a14284;
assign a18190 = a18188 & a14430;
assign a18192 = a18190 & a14288;
assign a18194 = a18192 & a14292;
assign a18196 = a18194 & a14310;
assign a18198 = a18196 & a14304;
assign a18200 = a18198 & a14298;
assign a18202 = a18200 & a14336;
assign a18204 = a18202 & a14372;
assign a18206 = a18204 & a14366;
assign a18208 = a18206 & a14360;
assign a18210 = a18208 & a14316;
assign a18212 = a18210 & a14320;
assign a18214 = a18212 & a14326;
assign a18216 = a18214 & a14332;
assign a18218 = a18216 & a14342;
assign a18220 = a18218 & a14348;
assign a18222 = a18220 & a14354;
assign a18224 = a18222 & a14378;
assign a18226 = a18224 & a14384;
assign a18228 = a18226 & a14390;
assign a18230 = a18228 & a14396;
assign a18232 = a18230 & a14402;
assign a18234 = a18232 & a14486;
assign a18236 = a18234 & a14448;
assign a18238 = a18236 & a14466;
assign a18240 = a18238 & a14408;
assign a18242 = a18240 & a14426;
assign a18244 = a18242 & a14420;
assign a18246 = a18244 & a14414;
assign a18248 = a18246 & a14242;
assign a18250 = a18170 & a17366;
assign a18252 = a18250 & a14238;
assign a18254 = a18252 & a14254;
assign a18256 = a18254 & a14248;
assign a18258 = a18256 & a14260;
assign a18260 = a18258 & a14266;
assign a18262 = a18260 & a14272;
assign a18264 = a18262 & a14278;
assign a18266 = a18264 & a14284;
assign a18268 = a18266 & a14430;
assign a18270 = a18268 & a14288;
assign a18272 = a18270 & a14292;
assign a18274 = a18272 & a14310;
assign a18276 = a18274 & a14304;
assign a18278 = a18276 & a14298;
assign a18280 = a18278 & a14336;
assign a18282 = a18280 & a14372;
assign a18284 = a18282 & a14366;
assign a18286 = a18284 & a14360;
assign a18288 = a18286 & a14316;
assign a18290 = a18288 & a14320;
assign a18292 = a18290 & a14326;
assign a18294 = a18292 & a14332;
assign a18296 = a18294 & a14342;
assign a18298 = a18296 & a14348;
assign a18300 = a18298 & a14354;
assign a18302 = a18300 & a14378;
assign a18304 = a18302 & a14384;
assign a18306 = a18304 & a14390;
assign a18308 = a18306 & a14396;
assign a18310 = a18308 & a14402;
assign a18312 = a18310 & a14486;
assign a18314 = a18312 & a14448;
assign a18316 = a18314 & a14466;
assign a18318 = a18316 & a14408;
assign a18320 = a18318 & a14426;
assign a18322 = a18320 & a14420;
assign a18324 = a18322 & a14414;
assign a18326 = a18324 & a14242;
assign a18328 = a18170 & a17450;
assign a18330 = a18328 & a14238;
assign a18332 = a18330 & a14254;
assign a18334 = a18332 & a14248;
assign a18336 = a18334 & a14260;
assign a18338 = a18336 & a14266;
assign a18340 = a18338 & a14272;
assign a18342 = a18340 & a14278;
assign a18344 = a18342 & a14284;
assign a18346 = a18344 & a14430;
assign a18348 = a18346 & a14288;
assign a18350 = a18348 & a14292;
assign a18352 = a18350 & a14310;
assign a18354 = a18352 & a14304;
assign a18356 = a18354 & a14298;
assign a18358 = a18356 & a14336;
assign a18360 = a18358 & a14372;
assign a18362 = a18360 & a14366;
assign a18364 = a18362 & a14360;
assign a18366 = a18364 & a14316;
assign a18368 = a18366 & a14320;
assign a18370 = a18368 & a14326;
assign a18372 = a18370 & a14332;
assign a18374 = a18372 & a14342;
assign a18376 = a18374 & a14348;
assign a18378 = a18376 & a14354;
assign a18380 = a18378 & a14378;
assign a18382 = a18380 & a14384;
assign a18384 = a18382 & a14390;
assign a18386 = a18384 & a14396;
assign a18388 = a18386 & a14402;
assign a18390 = a18388 & a14486;
assign a18392 = a18390 & a14448;
assign a18394 = a18392 & a14466;
assign a18396 = a18394 & a14408;
assign a18398 = a18396 & a14426;
assign a18400 = a18398 & a14420;
assign a18402 = a18400 & a14414;
assign a18404 = a18402 & a14242;
assign a18406 = a18170 & a17612;
assign a18408 = a18406 & a14238;
assign a18410 = a18408 & a14254;
assign a18412 = a18410 & a14248;
assign a18414 = a18412 & a14260;
assign a18416 = a18414 & a14266;
assign a18418 = a18416 & a14272;
assign a18420 = a18418 & a14278;
assign a18422 = a18420 & a14284;
assign a18424 = a18422 & a14430;
assign a18426 = a18424 & a14288;
assign a18428 = a18426 & a14292;
assign a18430 = a18428 & a14310;
assign a18432 = a18430 & a14304;
assign a18434 = a18432 & a14298;
assign a18436 = a18434 & a14336;
assign a18438 = a18436 & a14372;
assign a18440 = a18438 & a14366;
assign a18442 = a18440 & a14360;
assign a18444 = a18442 & a14316;
assign a18446 = a18444 & a14320;
assign a18448 = a18446 & a14326;
assign a18450 = a18448 & a14332;
assign a18452 = a18450 & a14342;
assign a18454 = a18452 & a14348;
assign a18456 = a18454 & a14354;
assign a18458 = a18456 & a14378;
assign a18460 = a18458 & a14384;
assign a18462 = a18460 & a14390;
assign a18464 = a18462 & a14396;
assign a18466 = a18464 & a14402;
assign a18468 = a18466 & a14486;
assign a18470 = a18468 & a14448;
assign a18472 = a18470 & a14466;
assign a18474 = a18472 & a14408;
assign a18476 = a18474 & a14426;
assign a18478 = a18476 & a14420;
assign a18480 = a18478 & a14414;
assign a18482 = a18480 & a14242;
assign a18484 = a18170 & a17852;
assign a18486 = a18484 & a14238;
assign a18488 = a18486 & a14254;
assign a18490 = a18488 & a14248;
assign a18492 = a18490 & a14260;
assign a18494 = a18492 & a14266;
assign a18496 = a18494 & a14272;
assign a18498 = a18496 & a14278;
assign a18500 = a18498 & a14284;
assign a18502 = a18500 & a14430;
assign a18504 = a18502 & a14288;
assign a18506 = a18504 & a14292;
assign a18508 = a18506 & a14310;
assign a18510 = a18508 & a14304;
assign a18512 = a18510 & a14298;
assign a18514 = a18512 & a14336;
assign a18516 = a18514 & a14372;
assign a18518 = a18516 & a14366;
assign a18520 = a18518 & a14360;
assign a18522 = a18520 & a14316;
assign a18524 = a18522 & a14320;
assign a18526 = a18524 & a14326;
assign a18528 = a18526 & a14332;
assign a18530 = a18528 & a14342;
assign a18532 = a18530 & a14348;
assign a18534 = a18532 & a14354;
assign a18536 = a18534 & a14378;
assign a18538 = a18536 & a14384;
assign a18540 = a18538 & a14390;
assign a18542 = a18540 & a14396;
assign a18544 = a18542 & a14402;
assign a18546 = a18544 & a14486;
assign a18548 = a18546 & a14448;
assign a18550 = a18548 & a14466;
assign a18552 = a18550 & a14408;
assign a18554 = a18552 & a14426;
assign a18556 = a18554 & a14420;
assign a18558 = a18556 & a14414;
assign a18560 = a18558 & a14242;
assign a18562 = ~a18560 & ~a18482;
assign a18564 = a18562 & ~a18404;
assign a18566 = a18564 & ~a18326;
assign a18568 = a18566 & ~a18248;
assign a18570 = a18568 & ~a18164;
assign a18572 = a18570 & ~a18086;
assign a18574 = a18572 & ~a18008;
assign a18576 = a18574 & ~a17930;
assign a18578 = a18576 & ~a17846;
assign a18580 = a18578 & ~a17768;
assign a18582 = a18580 & ~a17690;
assign a18584 = a18582 & ~a17606;
assign a18586 = a18584 & ~a17528;
assign a18588 = a18586 & ~a17444;
assign a18590 = a18588 & ~a17350;
assign a18592 = ~a18590 & a14214;
assign a18594 = ~l290 & ~i118;
assign a18596 = l290 & i118;
assign a18598 = ~a18596 & ~a18594;
assign a18600 = a14232 & a14226;
assign a18602 = a18600 & a14220;
assign a18604 = a18602 & a14254;
assign a18606 = a18604 & a14238;
assign a18608 = a18606 & a14248;
assign a18610 = a18608 & a14260;
assign a18612 = a18610 & a14266;
assign a18614 = a18612 & a14272;
assign a18616 = a18614 & a14278;
assign a18618 = a18616 & a14284;
assign a18620 = a18618 & a14430;
assign a18622 = a18620 & a14288;
assign a18624 = a18622 & a14292;
assign a18626 = a18624 & a14310;
assign a18628 = a18626 & a14304;
assign a18630 = a18628 & a14298;
assign a18632 = a18630 & a14336;
assign a18634 = a18632 & a14372;
assign a18636 = a18634 & a14366;
assign a18638 = a18636 & a14360;
assign a18640 = a18638 & a14316;
assign a18642 = a18640 & a14320;
assign a18644 = a18642 & a14326;
assign a18646 = a18644 & a14332;
assign a18648 = a18646 & a14342;
assign a18650 = a18648 & a14348;
assign a18652 = a18650 & a14354;
assign a18654 = a18652 & a14378;
assign a18656 = a18654 & a14384;
assign a18658 = a18656 & a14390;
assign a18660 = a18658 & a14396;
assign a18662 = a18660 & a14402;
assign a18664 = a18662 & a14486;
assign a18666 = a18664 & a14448;
assign a18668 = a18666 & a14466;
assign a18670 = a18668 & a14408;
assign a18672 = a18670 & a14426;
assign a18674 = a18672 & a14420;
assign a18676 = a18674 & a14414;
assign a18678 = a18676 & a14242;
assign a18680 = a18678 & a18598;
assign a18682 = ~a18680 & ~a18592;
assign a18684 = ~a18682 & a14208;
assign a18686 = ~l288 & ~i116;
assign a18688 = l288 & i116;
assign a18690 = ~a18688 & ~a18686;
assign a18692 = a14254 & a14214;
assign a18694 = a18692 & a14232;
assign a18696 = a18694 & a14226;
assign a18698 = a18696 & a14220;
assign a18700 = a18698 & a14238;
assign a18702 = a18700 & a14248;
assign a18704 = a18702 & a14260;
assign a18706 = a18704 & a14266;
assign a18708 = a18706 & a14272;
assign a18710 = a18708 & a14278;
assign a18712 = a18710 & a14284;
assign a18714 = a18712 & a14430;
assign a18716 = a18714 & a14288;
assign a18718 = a18716 & a14292;
assign a18720 = a18718 & a14310;
assign a18722 = a18720 & a14304;
assign a18724 = a18722 & a14298;
assign a18726 = a18724 & a14336;
assign a18728 = a18726 & a14372;
assign a18730 = a18728 & a14366;
assign a18732 = a18730 & a14360;
assign a18734 = a18732 & a14316;
assign a18736 = a18734 & a14320;
assign a18738 = a18736 & a14326;
assign a18740 = a18738 & a14332;
assign a18742 = a18740 & a14342;
assign a18744 = a18742 & a14348;
assign a18746 = a18744 & a14354;
assign a18748 = a18746 & a14378;
assign a18750 = a18748 & a14384;
assign a18752 = a18750 & a14390;
assign a18754 = a18752 & a14396;
assign a18756 = a18754 & a14402;
assign a18758 = a18756 & a14486;
assign a18760 = a18758 & a14448;
assign a18762 = a18760 & a14466;
assign a18764 = a18762 & a14408;
assign a18766 = a18764 & a14426;
assign a18768 = a18766 & a14420;
assign a18770 = a18768 & a14414;
assign a18772 = a18770 & a14242;
assign a18774 = a18772 & a18690;
assign a18776 = ~a18774 & ~a18684;
assign a18778 = ~a18776 & a14202;
assign a18780 = ~l238 & ~i66;
assign a18782 = l238 & i66;
assign a18784 = ~a18782 & ~a18780;
assign a18786 = a14214 & a14208;
assign a18788 = a18786 & a14254;
assign a18790 = a18788 & a14232;
assign a18792 = a18790 & a14226;
assign a18794 = a18792 & a14220;
assign a18796 = a18794 & a14238;
assign a18798 = a18796 & a14248;
assign a18800 = a18798 & a14260;
assign a18802 = a18800 & a14266;
assign a18804 = a18802 & a14272;
assign a18806 = a18804 & a14278;
assign a18808 = a18806 & a14284;
assign a18810 = a18808 & a14430;
assign a18812 = a18810 & a14288;
assign a18814 = a18812 & a14292;
assign a18816 = a18814 & a14310;
assign a18818 = a18816 & a14304;
assign a18820 = a18818 & a14298;
assign a18822 = a18820 & a14336;
assign a18824 = a18822 & a14372;
assign a18826 = a18824 & a14366;
assign a18828 = a18826 & a14360;
assign a18830 = a18828 & a14316;
assign a18832 = a18830 & a14320;
assign a18834 = a18832 & a14326;
assign a18836 = a18834 & a14332;
assign a18838 = a18836 & a14342;
assign a18840 = a18838 & a14348;
assign a18842 = a18840 & a14354;
assign a18844 = a18842 & a14378;
assign a18846 = a18844 & a14384;
assign a18848 = a18846 & a14390;
assign a18850 = a18848 & a14396;
assign a18852 = a18850 & a14402;
assign a18854 = a18852 & a14486;
assign a18856 = a18854 & a14448;
assign a18858 = a18856 & a14466;
assign a18860 = a18858 & a14408;
assign a18862 = a18860 & a14426;
assign a18864 = a18862 & a14420;
assign a18866 = a18864 & a14414;
assign a18868 = a18866 & a14242;
assign a18870 = a18868 & a18784;
assign a18872 = ~a18870 & ~a18778;
assign a18874 = ~a18872 & a14196;
assign a18876 = ~l216 & ~i44;
assign a18878 = l216 & i44;
assign a18880 = ~a18878 & ~a18876;
assign a18882 = a14208 & a14202;
assign a18884 = a18882 & a14214;
assign a18886 = a18884 & a14254;
assign a18888 = a18886 & a14232;
assign a18890 = a18888 & a14226;
assign a18892 = a18890 & a14220;
assign a18894 = a18892 & a14238;
assign a18896 = a18894 & a14248;
assign a18898 = a18896 & a14260;
assign a18900 = a18898 & a14266;
assign a18902 = a18900 & a14272;
assign a18904 = a18902 & a14278;
assign a18906 = a18904 & a14284;
assign a18908 = a18906 & a14430;
assign a18910 = a18908 & a14288;
assign a18912 = a18910 & a14292;
assign a18914 = a18912 & a14310;
assign a18916 = a18914 & a14304;
assign a18918 = a18916 & a14298;
assign a18920 = a18918 & a14336;
assign a18922 = a18920 & a14372;
assign a18924 = a18922 & a14366;
assign a18926 = a18924 & a14360;
assign a18928 = a18926 & a14316;
assign a18930 = a18928 & a14320;
assign a18932 = a18930 & a14326;
assign a18934 = a18932 & a14332;
assign a18936 = a18934 & a14342;
assign a18938 = a18936 & a14348;
assign a18940 = a18938 & a14354;
assign a18942 = a18940 & a14378;
assign a18944 = a18942 & a14384;
assign a18946 = a18944 & a14390;
assign a18948 = a18946 & a14396;
assign a18950 = a18948 & a14402;
assign a18952 = a18950 & a14486;
assign a18954 = a18952 & a14448;
assign a18956 = a18954 & a14466;
assign a18958 = a18956 & a14408;
assign a18960 = a18958 & a14426;
assign a18962 = a18960 & a14420;
assign a18964 = a18962 & a14414;
assign a18966 = a18964 & a14242;
assign a18968 = a18966 & a18880;
assign a18970 = ~a18968 & ~a18874;
assign a18972 = ~a18970 & a14190;
assign a18974 = ~l286 & ~i114;
assign a18976 = l286 & i114;
assign a18978 = ~a18976 & ~a18974;
assign a18980 = a14202 & a14196;
assign a18982 = a18980 & a14208;
assign a18984 = a18982 & a14214;
assign a18986 = a18984 & a14254;
assign a18988 = a18986 & a14232;
assign a18990 = a18988 & a14226;
assign a18992 = a18990 & a14220;
assign a18994 = a18992 & a14238;
assign a18996 = a18994 & a14248;
assign a18998 = a18996 & a14260;
assign a19000 = a18998 & a14266;
assign a19002 = a19000 & a14272;
assign a19004 = a19002 & a14278;
assign a19006 = a19004 & a14284;
assign a19008 = a19006 & a14430;
assign a19010 = a19008 & a14288;
assign a19012 = a19010 & a14292;
assign a19014 = a19012 & a14310;
assign a19016 = a19014 & a14304;
assign a19018 = a19016 & a14298;
assign a19020 = a19018 & a14336;
assign a19022 = a19020 & a14372;
assign a19024 = a19022 & a14366;
assign a19026 = a19024 & a14360;
assign a19028 = a19026 & a14316;
assign a19030 = a19028 & a14320;
assign a19032 = a19030 & a14326;
assign a19034 = a19032 & a14332;
assign a19036 = a19034 & a14342;
assign a19038 = a19036 & a14348;
assign a19040 = a19038 & a14354;
assign a19042 = a19040 & a14378;
assign a19044 = a19042 & a14384;
assign a19046 = a19044 & a14390;
assign a19048 = a19046 & a14396;
assign a19050 = a19048 & a14402;
assign a19052 = a19050 & a14486;
assign a19054 = a19052 & a14448;
assign a19056 = a19054 & a14466;
assign a19058 = a19056 & a14408;
assign a19060 = a19058 & a14426;
assign a19062 = a19060 & a14420;
assign a19064 = a19062 & a14414;
assign a19066 = a19064 & a14242;
assign a19068 = a19066 & a18978;
assign a19070 = ~a19068 & ~a18972;
assign a19072 = ~a19070 & a14184;
assign a19074 = ~l236 & ~i64;
assign a19076 = l236 & i64;
assign a19078 = ~a19076 & ~a19074;
assign a19080 = a14196 & a14190;
assign a19082 = a19080 & a14202;
assign a19084 = a19082 & a14208;
assign a19086 = a19084 & a14214;
assign a19088 = a19086 & a14254;
assign a19090 = a19088 & a14232;
assign a19092 = a19090 & a14226;
assign a19094 = a19092 & a14220;
assign a19096 = a19094 & a14238;
assign a19098 = a19096 & a14248;
assign a19100 = a19098 & a14260;
assign a19102 = a19100 & a14266;
assign a19104 = a19102 & a14272;
assign a19106 = a19104 & a14278;
assign a19108 = a19106 & a14284;
assign a19110 = a19108 & a14430;
assign a19112 = a19110 & a14288;
assign a19114 = a19112 & a14292;
assign a19116 = a19114 & a14310;
assign a19118 = a19116 & a14304;
assign a19120 = a19118 & a14298;
assign a19122 = a19120 & a14336;
assign a19124 = a19122 & a14372;
assign a19126 = a19124 & a14366;
assign a19128 = a19126 & a14360;
assign a19130 = a19128 & a14316;
assign a19132 = a19130 & a14320;
assign a19134 = a19132 & a14326;
assign a19136 = a19134 & a14332;
assign a19138 = a19136 & a14342;
assign a19140 = a19138 & a14348;
assign a19142 = a19140 & a14354;
assign a19144 = a19142 & a14378;
assign a19146 = a19144 & a14384;
assign a19148 = a19146 & a14390;
assign a19150 = a19148 & a14396;
assign a19152 = a19150 & a14402;
assign a19154 = a19152 & a14486;
assign a19156 = a19154 & a14448;
assign a19158 = a19156 & a14466;
assign a19160 = a19158 & a14408;
assign a19162 = a19160 & a14426;
assign a19164 = a19162 & a14420;
assign a19166 = a19164 & a14414;
assign a19168 = a19166 & a14242;
assign a19170 = a19168 & a19078;
assign a19172 = ~a19170 & ~a19072;
assign a19174 = ~a19172 & a14182;
assign a19176 = ~l284 & ~i112;
assign a19178 = l284 & i112;
assign a19180 = ~a19178 & ~a19176;
assign a19182 = a19180 & a14190;
assign a19184 = a19182 & a14184;
assign a19186 = a19184 & a14196;
assign a19188 = a19186 & a14202;
assign a19190 = a19188 & a14208;
assign a19192 = a19190 & a14214;
assign a19194 = a19192 & a14254;
assign a19196 = a19194 & a14232;
assign a19198 = a19196 & a14226;
assign a19200 = a19198 & a14220;
assign a19202 = a19200 & a14238;
assign a19204 = a19202 & a14248;
assign a19206 = a19204 & a14260;
assign a19208 = a19206 & a14266;
assign a19210 = a19208 & a14272;
assign a19212 = a19210 & a14278;
assign a19214 = a19212 & a14284;
assign a19216 = a19214 & a14430;
assign a19218 = a19216 & a14288;
assign a19220 = a19218 & a14292;
assign a19222 = a19220 & a14310;
assign a19224 = a19222 & a14304;
assign a19226 = a19224 & a14298;
assign a19228 = a19226 & a14336;
assign a19230 = a19228 & a14372;
assign a19232 = a19230 & a14366;
assign a19234 = a19232 & a14360;
assign a19236 = a19234 & a14316;
assign a19238 = a19236 & a14320;
assign a19240 = a19238 & a14326;
assign a19242 = a19240 & a14332;
assign a19244 = a19242 & a14342;
assign a19246 = a19244 & a14348;
assign a19248 = a19246 & a14354;
assign a19250 = a19248 & a14378;
assign a19252 = a19250 & a14384;
assign a19254 = a19252 & a14390;
assign a19256 = a19254 & a14396;
assign a19258 = a19256 & a14402;
assign a19260 = a19258 & a14486;
assign a19262 = a19260 & a14448;
assign a19264 = a19262 & a14466;
assign a19266 = a19264 & a14408;
assign a19268 = a19266 & a14426;
assign a19270 = a19268 & a14420;
assign a19272 = a19270 & a14414;
assign a19274 = a19272 & a14242;
assign a19276 = ~a19274 & ~a19174;
assign a19278 = ~l170 & l168;
assign a19280 = a19278 & l166;
assign a19282 = a19280 & ~l164;
assign a19284 = a19282 & ~a8022;
assign a19286 = a13108 & ~l166;
assign a19288 = a19286 & l164;
assign a19290 = a19288 & ~a8094;
assign a19292 = ~a19290 & ~a19284;
assign a19294 = ~a19292 & l172;
assign a19296 = ~a19294 & ~a19276;
assign a19298 = a14190 & a14184;
assign a19300 = a19298 & a14196;
assign a19302 = a19300 & a14202;
assign a19304 = a19302 & a14208;
assign a19306 = a19304 & a14214;
assign a19308 = a19306 & a14254;
assign a19310 = a19308 & a14232;
assign a19312 = a19310 & a14226;
assign a19314 = a19312 & a14220;
assign a19316 = a19314 & a14238;
assign a19318 = a19316 & a14248;
assign a19320 = a19318 & a14260;
assign a19322 = a19320 & a14266;
assign a19324 = a19322 & a14272;
assign a19326 = a19324 & a14278;
assign a19328 = a19326 & a14284;
assign a19330 = a19328 & a14430;
assign a19332 = a19330 & a14288;
assign a19334 = a19332 & a14292;
assign a19336 = a19334 & a14310;
assign a19338 = a19336 & a14304;
assign a19340 = a19338 & a14298;
assign a19342 = a19340 & a14336;
assign a19344 = a19342 & a14372;
assign a19346 = a19344 & a14366;
assign a19348 = a19346 & a14360;
assign a19350 = a19348 & a14316;
assign a19352 = a19350 & a14320;
assign a19354 = a19352 & a14326;
assign a19356 = a19354 & a14332;
assign a19358 = a19356 & a14342;
assign a19360 = a19358 & a14348;
assign a19362 = a19360 & a14354;
assign a19364 = a19362 & a14378;
assign a19366 = a19364 & a14384;
assign a19368 = a19366 & a14390;
assign a19370 = a19368 & a14396;
assign a19372 = a19370 & a14402;
assign a19374 = a19372 & a14486;
assign a19376 = a19374 & a14448;
assign a19378 = a19376 & a14466;
assign a19380 = a19378 & a14408;
assign a19382 = a19380 & a14426;
assign a19384 = a19382 & a14420;
assign a19386 = a19384 & a14414;
assign a19388 = a19386 & a14242;
assign a19390 = a19388 & a14182;
assign a19392 = a19390 & ~a19292;
assign a19394 = a19392 & l172;
assign a19396 = ~a19394 & ~a19296;
assign a19398 = ~a19396 & ~a14176;
assign a19400 = a19398 & ~a14174;
assign a19402 = a19400 & a14172;
assign a19404 = a19402 & a14160;
assign a19406 = a19404 & a14148;
assign a19408 = a19406 & a14138;
assign a19410 = a19408 & a14128;
assign a19412 = a19410 & a14116;
assign a19414 = a19412 & a14108;
assign a19416 = a19414 & a14100;
assign a19418 = a19416 & a14090;
assign a19420 = a19418 & a14080;
assign a19422 = a19420 & ~a698;
assign a19424 = a19422 & ~a696;
assign a19426 = a19424 & a14070;
assign a19428 = a19426 & a14052;
assign a19430 = a19428 & a14036;
assign a19432 = a19430 & a14000;
assign a19434 = a19432 & a13962;
assign a19436 = a19434 & a13940;
assign a19438 = a19436 & a13914;
assign a19440 = a19438 & a13892;
assign a19442 = a19440 & a13782;
assign a19444 = a19442 & a13088;
assign a19446 = a19444 & a12404;
assign a19448 = a19446 & a11640;
assign a19450 = a19448 & a10640;
assign a19452 = a19450 & a7856;
assign a19454 = a19452 & a7602;
assign a19456 = a19454 & a7364;
assign a19458 = a19456 & a6654;
assign a19460 = a19458 & a5882;
assign a19462 = a19460 & a5048;
assign a19464 = a19462 & a4288;
assign a19466 = a19464 & a3308;
assign a19468 = a19466 & l338;
assign a19470 = ~a19468 & l340;
assign a19474 = ~l274 & ~l272;
assign a19476 = a2384 & a2304;
assign a19478 = a19476 & a2520;
assign a19480 = a19478 & a2682;
assign a19482 = a19480 & a4346;
assign a19484 = a19482 & a850;
assign a19486 = a19484 & a1004;
assign a19488 = a19486 & a1070;
assign a19490 = a19488 & a1206;
assign a19492 = a19490 & a1450;
assign a19494 = a19492 & a1514;
assign a19496 = a19494 & a1652;
assign a19498 = a19496 & a1774;
assign a19500 = a19498 & a1898;
assign a19502 = a19500 & a1990;
assign a19504 = a19502 & a2060;
assign a19506 = a19504 & a6030;
assign a19508 = ~a19506 & a19474;
assign a19510 = a2384 & a2236;
assign a19512 = a19510 & a2520;
assign a19514 = a19512 & a2682;
assign a19516 = a19514 & a4346;
assign a19518 = a19516 & a850;
assign a19520 = a19518 & a1004;
assign a19522 = a19520 & a1070;
assign a19524 = a19522 & a1206;
assign a19526 = a19524 & a1450;
assign a19528 = a19526 & a1514;
assign a19530 = a19528 & a1652;
assign a19532 = a19530 & a1774;
assign a19534 = a19532 & a1898;
assign a19536 = a19534 & a1990;
assign a19538 = a19536 & a2060;
assign a19540 = a19538 & a6030;
assign a19542 = l274 & l272;
assign a19544 = a19542 & ~a19540;
assign a19546 = ~a19544 & ~a19508;
assign a19548 = ~a19546 & l276;
assign a19550 = a2306 & a2236;
assign a19552 = a19550 & a2520;
assign a19554 = a19552 & a2682;
assign a19556 = a19554 & a4346;
assign a19558 = a19556 & a850;
assign a19560 = a19558 & a1004;
assign a19562 = a19560 & a1070;
assign a19564 = a19562 & a1206;
assign a19566 = a19564 & a1450;
assign a19568 = a19566 & a1514;
assign a19570 = a19568 & a1652;
assign a19572 = a19570 & a1774;
assign a19574 = a19572 & a1898;
assign a19576 = a19574 & a1990;
assign a19578 = a19576 & a2060;
assign a19580 = a19578 & a6030;
assign a19582 = ~a19580 & a846;
assign a19584 = a19550 & a2384;
assign a19586 = a19584 & a2682;
assign a19588 = a19586 & a4346;
assign a19590 = a19588 & a850;
assign a19592 = a19590 & a1004;
assign a19594 = a19592 & a1070;
assign a19596 = a19594 & a1206;
assign a19598 = a19596 & a1450;
assign a19600 = a19598 & a1514;
assign a19602 = a19600 & a1652;
assign a19604 = a19602 & a1774;
assign a19606 = a19604 & a1898;
assign a19608 = a19606 & a1990;
assign a19610 = a19608 & a2060;
assign a19612 = a19610 & a6030;
assign a19614 = ~a19612 & a1202;
assign a19616 = ~a19614 & ~a19582;
assign a19618 = a19616 & ~a19548;
assign a19620 = ~a19618 & l270;
assign a19622 = a19620 & ~l268;
assign a19624 = a19584 & a2520;
assign a19626 = a19624 & a4346;
assign a19628 = a19626 & a850;
assign a19630 = a19628 & a1004;
assign a19632 = a19630 & a1070;
assign a19634 = a19632 & a1206;
assign a19636 = a19634 & a1450;
assign a19638 = a19636 & a1514;
assign a19640 = a19638 & a1652;
assign a19642 = a19640 & a1774;
assign a19644 = a19642 & a1898;
assign a19646 = a19644 & a1990;
assign a19648 = a19646 & a2060;
assign a19650 = a19648 & a6030;
assign a19652 = ~a19650 & a2682;
assign a19654 = a19624 & a2682;
assign a19656 = a19654 & a850;
assign a19658 = a19656 & a1004;
assign a19660 = a19658 & a1070;
assign a19662 = a19660 & a1206;
assign a19664 = a19662 & a1450;
assign a19666 = a19664 & a1514;
assign a19668 = a19666 & a1652;
assign a19670 = a19668 & a1774;
assign a19672 = a19670 & a1898;
assign a19674 = a19672 & a1990;
assign a19676 = a19674 & a2060;
assign a19678 = a19676 & a6030;
assign a19680 = ~a19678 & a4346;
assign a19682 = a19654 & a4346;
assign a19684 = a19682 & a1004;
assign a19686 = a19684 & a1070;
assign a19688 = a19686 & a1206;
assign a19690 = a19688 & a1450;
assign a19692 = a19690 & a1514;
assign a19694 = a19692 & a1652;
assign a19696 = a19694 & a1774;
assign a19698 = a19696 & a1898;
assign a19700 = a19698 & a1990;
assign a19702 = a19700 & a2060;
assign a19704 = a19702 & a6030;
assign a19706 = ~a19704 & a850;
assign a19708 = a19682 & a850;
assign a19710 = a19708 & a1070;
assign a19712 = a19710 & a1206;
assign a19714 = a19712 & a1450;
assign a19716 = a19714 & a1514;
assign a19718 = a19716 & a1652;
assign a19720 = a19718 & a1774;
assign a19722 = a19720 & a1898;
assign a19724 = a19722 & a1990;
assign a19726 = a19724 & a2060;
assign a19728 = a19726 & a6030;
assign a19730 = ~a19728 & a1004;
assign a19732 = a19708 & a1004;
assign a19734 = a19732 & a1206;
assign a19736 = a19734 & a1450;
assign a19738 = a19736 & a1514;
assign a19740 = a19738 & a1652;
assign a19742 = a19740 & a1774;
assign a19744 = a19742 & a1898;
assign a19746 = a19744 & a1990;
assign a19748 = a19746 & a2060;
assign a19750 = a19748 & a6030;
assign a19752 = ~a19750 & a1070;
assign a19754 = a19732 & a1070;
assign a19756 = a19754 & a1450;
assign a19758 = a19756 & a1514;
assign a19760 = a19758 & a1652;
assign a19762 = a19760 & a1774;
assign a19764 = a19762 & a1898;
assign a19766 = a19764 & a1990;
assign a19768 = a19766 & a2060;
assign a19770 = a19768 & a6030;
assign a19772 = ~a19770 & a1206;
assign a19774 = a19754 & a1206;
assign a19776 = a19774 & a1514;
assign a19778 = a19776 & a1652;
assign a19780 = a19778 & a1774;
assign a19782 = a19780 & a1898;
assign a19784 = a19782 & a1990;
assign a19786 = a19784 & a2060;
assign a19788 = a19786 & a6030;
assign a19790 = ~a19788 & a1450;
assign a19792 = a19774 & a1450;
assign a19794 = a19792 & a1652;
assign a19796 = a19794 & a1774;
assign a19798 = a19796 & a1898;
assign a19800 = a19798 & a1990;
assign a19802 = a19800 & a2060;
assign a19804 = a19802 & a6030;
assign a19806 = ~a19804 & a1514;
assign a19808 = a19792 & a1514;
assign a19810 = a19808 & a1774;
assign a19812 = a19810 & a1898;
assign a19814 = a19812 & a1990;
assign a19816 = a19814 & a2060;
assign a19818 = a19816 & a6030;
assign a19820 = ~a19818 & a1652;
assign a19822 = a19808 & a1652;
assign a19824 = a19822 & a1898;
assign a19826 = a19824 & a1990;
assign a19828 = a19826 & a2060;
assign a19830 = a19828 & a6030;
assign a19832 = ~a19830 & a1774;
assign a19834 = a19822 & a1774;
assign a19836 = a19834 & a1990;
assign a19838 = a19836 & a2060;
assign a19840 = a19838 & a6030;
assign a19842 = ~a19840 & a1898;
assign a19844 = a19834 & a1898;
assign a19846 = a19844 & a2060;
assign a19848 = a19846 & a6030;
assign a19850 = ~a19848 & a1990;
assign a19852 = a19844 & a1990;
assign a19854 = a19852 & a6030;
assign a19856 = ~a19854 & a2060;
assign a19858 = a19852 & a2060;
assign a19860 = ~a19858 & a6030;
assign a19862 = ~a19860 & ~a19856;
assign a19864 = a19862 & ~a19850;
assign a19866 = a19864 & ~a19842;
assign a19868 = a19866 & ~a19832;
assign a19870 = a19868 & ~a19820;
assign a19872 = a19870 & ~a19806;
assign a19874 = a19872 & ~a19790;
assign a19876 = a19874 & ~a19772;
assign a19878 = a19876 & ~a19752;
assign a19880 = a19878 & ~a19730;
assign a19882 = a19880 & ~a19706;
assign a19884 = a19882 & ~a19680;
assign a19886 = a19884 & ~a19652;
assign a19888 = a19886 & ~a19622;
assign a19890 = a19888 & l338;
assign a19892 = ~a13108 & ~a7860;
assign a19894 = ~a19892 & l166;
assign a19896 = a19894 & ~l164;
assign a19898 = l250 & l248;
assign a19900 = ~a19898 & ~a7626;
assign a19902 = a19900 & ~l252;
assign a19904 = ~a19902 & ~a7108;
assign a19906 = a19904 & ~a7146;
assign a19908 = a19906 & ~a7018;
assign a19910 = ~a19908 & ~a19896;
assign a19912 = a19910 & ~a9354;
assign a19914 = a19912 & ~a6726;
assign a19916 = a19914 & ~a9458;
assign a19918 = a19916 & ~a8776;
assign a19920 = a19918 & ~a9556;
assign a19922 = a19920 & ~a8846;
assign a19924 = a19922 & ~a9636;
assign a19926 = a19924 & ~a8932;
assign a19928 = a19926 & ~a11688;
assign a19930 = a19928 & ~a9154;
assign a19932 = a19930 & ~a8998;
assign a19934 = a19932 & ~a9070;
assign a19936 = a19908 & a8550;
assign a19938 = a19908 & a11728;
assign a19940 = a19908 & a8626;
assign a19942 = a19908 & a9354;
assign a19944 = a19908 & a6726;
assign a19946 = a19908 & a9556;
assign a19948 = a19908 & a9458;
assign a19950 = a19908 & a8776;
assign a19952 = a19908 & a8846;
assign a19954 = a19908 & a9636;
assign a19956 = a19908 & a8932;
assign a19958 = a19908 & a11688;
assign a19960 = a19908 & a9154;
assign a19962 = a19908 & a8998;
assign a19964 = a19908 & a9070;
assign a19966 = a19908 & ~a8550;
assign a19968 = a19966 & ~a11728;
assign a19970 = a19968 & ~a8626;
assign a19972 = a19970 & ~a9354;
assign a19974 = a19972 & ~a6726;
assign a19976 = a19974 & ~a9458;
assign a19978 = a19976 & ~a8776;
assign a19980 = a19978 & ~a9556;
assign a19982 = a19980 & ~a8846;
assign a19984 = a19982 & ~a9636;
assign a19986 = a19984 & ~a8932;
assign a19988 = a19986 & ~a11688;
assign a19990 = a19988 & ~a9154;
assign a19992 = a19990 & ~a8998;
assign a19994 = a19992 & ~a9070;
assign a19996 = ~a19994 & ~a19964;
assign a19998 = a19996 & ~a19962;
assign a20000 = a19998 & ~a19960;
assign a20002 = a20000 & ~a19958;
assign a20004 = a20002 & ~a19956;
assign a20006 = a20004 & ~a19954;
assign a20008 = a20006 & ~a19952;
assign a20010 = a20008 & ~a19950;
assign a20012 = a20010 & ~a19948;
assign a20014 = a20012 & ~a19946;
assign a20016 = a20014 & ~a19944;
assign a20018 = a20016 & ~a19942;
assign a20020 = a20018 & ~a19940;
assign a20022 = a20020 & ~a19938;
assign a20024 = a20022 & ~a19936;
assign a20026 = a20024 & ~a19934;
assign a20028 = a20026 & l338;
assign a20030 = l170 & ~l164;
assign a20032 = l172 & ~l168;
assign a20034 = a20032 & ~l166;
assign a20036 = ~l172 & l168;
assign a20038 = a20036 & l166;
assign a20040 = ~a20038 & ~a20034;
assign a20042 = ~a20040 & a20030;
assign a20044 = ~a20042 & a7060;
assign a20046 = a20044 & l338;
assign a20048 = a9244 & a9184;
assign a20050 = a20048 & l338;
assign a20052 = ~a19278 & ~a6722;
assign a20054 = a20052 & ~a9150;
assign a20056 = a20054 & ~a9240;
assign a20058 = a20056 & ~a9066;
assign a20060 = ~a20058 & l166;
assign a20062 = ~a20060 & ~a8996;
assign a20064 = a20062 & ~a8930;
assign a20066 = a20064 & ~a8844;
assign a20068 = a20066 & ~a7862;
assign a20070 = a20068 & ~a6724;
assign a20072 = a20070 & ~a9152;
assign a20074 = a20072 & ~a9302;
assign a20076 = a20074 & ~a9184;
assign a20078 = ~a20064 & ~l164;
assign a20080 = a20078 & ~a8844;
assign a20082 = a20080 & ~a8776;
assign a20084 = a20082 & ~a6726;
assign a20086 = a20084 & ~a9154;
assign a20088 = a20086 & ~a9304;
assign a20090 = a20088 & ~a9186;
assign a20092 = ~a13094 & ~a9636;
assign a20094 = a20092 & ~a9556;
assign a20096 = ~a20094 & ~a8010;
assign a20098 = a20096 & ~a8626;
assign a20100 = a20098 & ~a8550;
assign a20102 = a20100 & ~a11728;
assign a20104 = ~a20102 & ~a9244;
assign a20106 = a20104 & ~a9070;
assign a20108 = a20106 & ~a8998;
assign a20110 = a20108 & ~a8932;
assign a20112 = ~a20110 & ~a8846;
assign a20114 = a20112 & ~a8776;
assign a20116 = a20114 & ~a6726;
assign a20118 = a20116 & ~a9154;
assign a20120 = ~a20118 & ~a9304;
assign a20122 = a20034 & ~l164;
assign a20124 = l172 & l168;
assign a20126 = a20124 & ~l166;
assign a20128 = a20126 & ~l164;
assign a20130 = a20032 & l166;
assign a20132 = a20130 & ~l164;
assign a20134 = a20124 & l166;
assign a20136 = a20134 & ~l164;
assign a20138 = ~l168 & ~l166;
assign a20140 = a20138 & l164;
assign a20142 = a20140 & ~a9302;
assign a20144 = a20142 & ~a11688;
assign a20146 = a20038 & ~l164;
assign a20148 = ~a20146 & ~a20144;
assign a20150 = a20148 & ~a20136;
assign a20152 = ~a20150 & ~a8010;
assign a20154 = a20152 & ~a8626;
assign a20156 = a9712 & l166;
assign a20158 = a20156 & ~l164;
assign a20160 = ~a20158 & ~a20154;
assign a20162 = a20160 & ~a20132;
assign a20164 = ~a20162 & ~a9244;
assign a20166 = a20164 & ~a9070;
assign a20168 = a20036 & ~l166;
assign a20170 = a20168 & ~l164;
assign a20172 = ~a20170 & ~a20166;
assign a20174 = a20172 & ~a20128;
assign a20176 = ~a20174 & ~a8846;
assign a20178 = a20176 & ~a8776;
assign a20180 = a9712 & ~l166;
assign a20182 = a20180 & ~l164;
assign a20184 = ~a20182 & ~a20178;
assign a20186 = a20184 & ~a20122;
assign a20188 = a13092 & ~l164;
assign a20190 = a19286 & ~l164;
assign a20192 = a19278 & ~l166;
assign a20194 = a20192 & ~l164;
assign a20196 = l170 & l168;
assign a20198 = a20196 & ~l166;
assign a20200 = a20198 & ~l164;
assign a20202 = a13090 & l166;
assign a20204 = a20202 & ~l164;
assign a20206 = a20196 & l166;
assign a20208 = a20206 & ~l164;
assign a20210 = a9458 & l170;
assign a20212 = ~a20210 & a20140;
assign a20214 = a20212 & ~a11688;
assign a20216 = ~a20214 & ~a20208;
assign a20218 = ~a20216 & ~a9556;
assign a20220 = ~a20218 & ~a19282;
assign a20222 = ~a20220 & ~a8626;
assign a20224 = ~a20222 & ~a13112;
assign a20226 = ~a20224 & ~a11728;
assign a20228 = ~a20226 & ~a20204;
assign a20230 = ~a20228 & ~a9070;
assign a20232 = ~a20230 & ~a20200;
assign a20234 = ~a20232 & ~a8932;
assign a20236 = ~a20234 & ~a20194;
assign a20238 = ~a20236 & ~a8776;
assign a20240 = ~a20238 & ~a20190;
assign a20242 = ~a20240 & ~a9154;
assign a20244 = ~a20242 & ~a20188;
assign a20246 = ~a20244 & l172;
assign a20248 = a20246 & ~a9186;
assign a20250 = ~a20248 & ~l204;
assign a20252 = a20248 & l204;
assign a20254 = ~a20252 & ~a20250;
assign a20256 = ~a20254 & ~a20186;
assign a20258 = a20256 & l170;
assign a20260 = a20258 & ~a9304;
assign a20262 = a20260 & ~a9186;
assign a20264 = a20262 & ~a20120;
assign a20266 = a20264 & ~a20090;
assign a20268 = a20266 & ~a20076;
assign a20270 = a20268 & ~l164;
assign a20272 = ~a20270 & ~a20042;
assign a20274 = a20272 & ~a9354;
assign a20276 = a20274 & ~a9458;
assign a20278 = a20276 & ~a8550;
assign a20280 = a20278 & ~a8626;
assign a20282 = a20280 & ~a8776;
assign a20284 = a20282 & ~a9636;
assign a20286 = a20284 & ~a8998;
assign a20288 = a20286 & ~a9070;
assign a20290 = a20288 & ~a8846;
assign a20292 = a20290 & ~a11688;
assign a20294 = a20292 & ~a8932;
assign a20296 = l276 & ~l270;
assign a20298 = ~l276 & l270;
assign a20300 = ~a20298 & ~a20296;
assign a20302 = ~a20300 & ~l272;
assign a20304 = ~a20302 & ~a5094;
assign a20306 = ~a20304 & l274;
assign a20308 = a20306 & ~l268;
assign a20310 = a20308 & ~a20294;
assign a20312 = a20310 & l338;
assign a20314 = ~a7858 & l168;
assign a20316 = ~a20314 & ~l166;
assign a20318 = ~a20316 & l164;
assign a20320 = ~l182 & ~l180;
assign a20322 = ~a20320 & l178;
assign a20324 = ~a20322 & ~l176;
assign a20326 = ~a20324 & l174;
assign a20328 = a14092 & l188;
assign a20330 = a7948 & l242;
assign a20332 = a7106 & l248;
assign a20334 = ~a6728 & l254;
assign a20336 = a19474 & ~l270;
assign a20338 = ~a20336 & l268;
assign a20340 = l280 & l278;
assign a20342 = ~a20340 & ~a20338;
assign a20344 = a20342 & ~a20334;
assign a20346 = a20344 & ~a20332;
assign a20348 = a20346 & ~a20330;
assign a20350 = a20348 & ~a20328;
assign a20352 = a20350 & ~a20326;
assign a20354 = a20352 & ~a20318;
assign a20356 = ~a20354 & l340;
assign p0 = a19890;
assign p1 = a20028;
assign p2 = a20046;
assign p3 = a20050;
assign p4 = a20312;

assert property (~p0);
assert property (~p1);
assert property (~p2);
assert property (~p3);
assert property (~p4);

endmodule
