module main;

  typedef bit some_identifier;

  // name collision
  typedef bit some_identifier;

endmodule
