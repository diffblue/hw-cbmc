module main();

   // IEEE 1800-2017 A.2.2.1
   shortreal some_shortreal;
   real some_real;
   realtime some_realtime;

endmodule
