module main;
  // The empty item.
  ;

  generate
    // Also inside generate
    ;
  endgenerate

endmodule
