module my_module(input x, y);

endmodule

module main();

  my_module m(1);

endmodule
