module main;

  typedef enum { some_identifier } some_type;

  // name collision
  wire some_identifier;

endmodule
