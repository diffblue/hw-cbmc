module main;

  // powers with constant rhs
  property1: assert final (3**0==1);
  property2: assert final (3**1==3);
  property3: assert final ((-3)**1==-3);
  property4: assert final (3**3==27);

endmodule
