package some_package;

typedef int some_type;

typedef struct packed {
  some_type some_field;
} other_type;

endpackage

module top;
endmodule
