module top;
  sub instance1();
  sub instance2();
endmodule

module sub;
  subsub instance3();
endmodule 

module subsub;
endmodule
