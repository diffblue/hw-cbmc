module main(input clk);

  initial p0: assert property (s_nexttime 0);

endmodule
