module some_module;
  // endmodule identifiers are a SystemVerilog feature
endmodule : some_module

