module top;
  import my_package::*;
  my_package::some_type some_var;
endmodule
