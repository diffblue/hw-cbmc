module main;

  // 1800-2017 6.12.1
  real some_real;
  wire [7:0] x = some_real[7:0];

endmodule
