module main;

  int string_to_int[string]; 
  string integral_to_string[*];

endmodule
