module top;
  interconnect bus;
  mod1 m1(bus);
  mod2 m2(bus);
endmodule

module mod1(input in);
endmodule

module mod2(output out);
endmodule
