// default values for inputs must be constants
module M(input a, input b = a);

endmodule
