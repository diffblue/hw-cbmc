module main;
  assert property ({5'bxz01?, 4'b10zx} === 9'bxz01?10zx);
endmodule
