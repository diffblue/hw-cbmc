module main;

  parameter p = 123;
  parameter p = 123;

endmodule
