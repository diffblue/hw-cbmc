module main;

  initial $display("Internal error: null handle at %s, line %d.",
    `__FILE__, `__LINE__);

endmodule
