module bobmiterbm1multi (i2,i4,i6,i8,i10,i12,i14,i16,i18,i20,i22,i24,i26,i28,i30,
i32,i34,i36,i38,i40,i42,i44,i46,i48,i50,i52,i54,i56,i58,i60,
i62,i64,i66,i68,i70,i72,i74,i76,i78,i80,i82,i84,i86,i88,i90,
i92,i94,i96,i98,i100,i102,i104,i106,i108,i110,i112,i114,i116,i118,i120,
i122,i124,i126,i128,i130,i132,i134,i136,i138,i140,i142,i144,i146,i148,i150,
i152,i154,i156,i158,i160,i162,i164,i166,i168,i170,i172,i174,i176,i178,i180,
i182,i184,i186,i188,i190,i192,i194,i196,i198,i200,i202,i204,i206,i208,i210,
i212,i214,i216,i218,i220,i222,i224,i226,i228,i230,i232,i234,i236,i238,i240,
i242,i244,p0,p1,p2,p3,p4,p5,p6,p7,p8,p9,p10,p11,p12,
p13,p14,p15,p16,p17,p18,p19,p20,p21,p22,p23,p24,p25,p26,p27,
p28,p29,p30,p31,p32,p33,p34,p35,p36,p37,p38,p39,p40,p41,p42,
p43,p44,p45,p46,p47,p48,p49,p50,p51,p52,p53,p54,p55,p56,p57,
p58,p59,p60,p61,p62,p63,p64,p65,p66,p67,p68,p69,p70,p71,p72,
p73,p74,p75,p76,p77,p78,p79,p80,p81,p82,p83,p84,p85,p86,p87,
p88,p89,p90,p91,p92,p93,p94,p95,p96,p97,p98,p99,p100,p101,p102,
p103,p104,p105,p106,p107,p108,p109,p110,p111,p112,p113,p114,p115,p116,p117,
p118,p119,p120,p121,p122,p123,p124,p125,p126,p127,p128,p129,p130,p131,p132,
p133,p134,p135,p136,p137,p138,p139,p140,p141,p142,p143,p144,p145,p146,p147,
p148,p149,p150,p151,p152,p153,p154,p155,p156,p157,p158,p159,p160,p161,p162,
p163,p164,p165,p166,p167,p168,p169,p170,p171,p172,p173,p174,p175,p176,p177,
p178,p179,p180,p181,p182,p183,p184,p185,p186,p187,p188,p189,p190,p191,p192,
p193,p194,p195,p196,p197,p198,p199,p200,p201,p202,p203,p204,p205,p206,p207,
p208,p209,p210,p211,p212,p213,p214,p215,p216,p217,p218,p219,p220,p221,p222,
p223,p224,p225,p226,p227,p228,p229,p230,p231,p232,p233,p234,p235,p236,p237,
p238,p239,p240,p241,p242,p243,p244,p245,p246,p247,p248,p249,p250,p251,p252,
p253,p254,p255,p256,p257,p258,p259,p260,p261,p262,p263,p264,p265,p266,p267,
p268,p269,p270,p271,p272,p273,p274,p275,p276,p277,p278,p279,p280,p281,p282,
p283,p284,p285,p286,p287,p288,p289,p290,p291,p292,p293,p294,p295,p296,p297,
p298,p299,p300,p301,p302,p303,p304,p305,p306,p307,p308,p309,p310,p311,p312,
p313,p314,p315,p316,p317,p318,p319,p320,p321,p322,p323,p324,p325,p326,p327,
p328,p329,p330,p331,p332,p333,p334,p335,p336,p337,p338,p339,p340,p341,p342,
p343,p344,p345,p346,p347,p348,p349,p350,p351,p352,p353,p354,p355,p356,p357,
p358,p359,p360,p361,p362,p363,p364,p365,p366,p367,p368,p369,p370,p371,p372,
p373,p374,p375,p376,p377,p378,p379,p380,p381,p382,p383,p384,p385,p386,p387,
p388,p389,p390,p391,p392,p393,p394,p395,p396,p397,p398,p399,p400,p401,p402,
p403,p404,p405,p406,p407,p408,p409,p410,p411,p412,p413,p414,p415,p416,p417,
p418,p419,p420,p421,p422,p423,p424,p425,p426,p427,p428,p429,p430,p431,p432,
p433,p434,p435,p436,p437,p438,p439,p440,p441,p442,p443,p444,p445,p446,p447,
p448,p449,p450,p451,p452,p453,p454,p455,p456,p457,p458,p459,p460,p461,p462,
p463,p464,p465,p466,p467,p468,p469,p470,p471,p472,p473,p474,p475,p476,p477,
p478,p479,p480,p481,p482,p483,p484,p485,p486,p487,p488,p489,p490,p491,p492,
p493,p494,p495,p496,p497,p498,p499,p500,p501,p502,p503,p504,p505,p506,p507,
p508,p509,p510,p511,p512,p513,p514,p515,p516,p517,p518,p519,p520,p521,p522,
p523,p524,p525,p526,p527,p528,p529,p530,p531,p532,p533,p534,p535,p536,p537,
p538,p539,p540,p541,p542,p543,p544,p545,p546,p547,p548,p549,p550,p551,p552,
p553,p554,p555,p556,p557,p558,p559,p560,p561,p562,p563,p564,p565,p566,p567,
p568,p569,p570,p571,p572,p573,p574,p575,p576,p577,p578,p579,p580,p581,p582,
p583,p584,p585,p586,p587,p588,p589,p590,p591,p592,p593,p594,p595,p596,p597,
p598,p599,p600,p601,p602,p603,p604,p605,p606,p607,p608,p609,p610,p611,p612,
p613,p614,p615,p616,p617,p618,p619,p620,p621,p622,p623,p624,p625,p626,p627,
p628,p629,p630,p631,p632,p633,p634,p635,p636,p637,p638,p639,p640,p641,p642,
p643,p644,p645,p646,p647,p648,p649,p650,p651,p652,p653,p654,p655,p656,p657,
p658,p659,p660,p661,p662,p663,p664,p665,p666,p667,p668,p669,p670,p671,p672,
p673,p674,p675,p676,p677,p678,p679,p680,p681,p682,p683,p684,p685,p686,p687,
p688,p689,p690,p691,p692,p693,p694,p695,p696,p697,p698,p699,p700,p701,p702,
p703,p704,p705,p706,p707,p708,p709,p710,p711,p712,p713,p714,p715,p716,p717,
p718,p719,p720,p721,p722,p723,p724,p725,p726,p727,p728,p729,p730,p731,p732,
p733,p734,p735,p736,p737,p738,p739,p740,p741,p742,p743,p744,p745,p746,p747,
p748,p749,p750,p751,p752,p753,p754,p755,p756,p757,p758,p759,p760,p761,p762,
p763,p764,p765,p766,p767,p768,p769,p770,p771,p772,p773,p774,p775,p776,p777,
p778,p779,p780,p781,p782,p783,p784,p785,p786,p787,p788,p789,p790,p791,p792,
p793,p794,p795,p796,p797,p798,p799,p800,p801,p802,p803,p804,p805,p806,p807,
p808,p809,p810,p811,p812,p813,p814,p815,p816,p817,p818,p819,p820,p821,p822,
p823,p824,p825,p826,p827,p828,p829,p830,p831,p832,p833,p834,p835,p836,p837,
p838,p839,p840,p841,p842,p843,p844,p845,p846,p847,p848,p849,p850,p851,p852,
p853,p854,p855,p856,p857,p858,p859,p860,p861,p862,p863,p864,p865,p866,p867,
p868,p869,p870,p871,p872,p873,p874,p875,p876,p877,p878,p879,p880,p881,p882,
p883,p884,p885,p886,p887,p888,p889,p890,p891,p892,p893,p894,p895,p896,p897,
p898,p899,p900,p901,p902,p903,p904,p905,p906,p907,p908,p909,p910,p911,p912,
p913,p914,p915,p916,p917,p918,p919,p920,p921,p922,p923,p924,p925,p926,p927,
p928,p929,p930,p931,p932,p933,p934,p935,p936,p937,p938,p939,p940,p941,p942,
p943,p944,p945,p946,p947,p948,p949,p950,p951,p952,p953,p954,p955,p956,p957,
p958,p959,p960,p961,p962,p963,p964,p965,p966,p967,p968,p969,p970,p971,p972,
p973,p974,p975,p976,p977,p978,p979,p980,p981,p982,p983,p984,p985,p986,p987,
p988,p989,p990,p991,p992,p993,p994,p995,p996,p997,p998,p999,p1000,p1001,p1002,
p1003,p1004,p1005,p1006,p1007,p1008,p1009,p1010,p1011,p1012,p1013,p1014,p1015,p1016,p1017,
p1018,p1019,p1020,p1021,p1022,p1023,p1024,p1025,p1026,p1027,p1028,p1029,p1030,p1031,p1032,
p1033,p1034,p1035,p1036,p1037,p1038,p1039,p1040,p1041,p1042,p1043,p1044,p1045,p1046,p1047,
p1048,p1049,p1050,p1051,p1052,p1053,p1054,p1055,p1056,p1057,p1058,p1059,p1060,p1061,p1062,
p1063,p1064,p1065,p1066,p1067,p1068,p1069,p1070,p1071,p1072,p1073,p1074,p1075,p1076,p1077,
p1078,p1079,p1080,p1081,p1082,p1083,p1084,p1085,p1086,p1087,p1088,p1089,p1090,p1091,p1092,
p1093,p1094,p1095,p1096,p1097,p1098,p1099,p1100,p1101,p1102,p1103,p1104,p1105,p1106,p1107,
p1108,p1109,p1110,p1111,p1112,p1113,p1114,p1115,p1116,p1117,p1118,p1119,p1120,p1121,p1122,
p1123,p1124,p1125,p1126,p1127,p1128,p1129,p1130,p1131,p1132,p1133,p1134,p1135,p1136,p1137,
p1138,p1139,p1140,p1141,p1142,p1143,p1144,p1145,p1146,p1147,p1148,p1149);

input i2,i4,i6,i8,i10,i12,i14,i16,i18,i20,i22,i24,i26,i28,i30,
i32,i34,i36,i38,i40,i42,i44,i46,i48,i50,i52,i54,i56,i58,i60,
i62,i64,i66,i68,i70,i72,i74,i76,i78,i80,i82,i84,i86,i88,i90,
i92,i94,i96,i98,i100,i102,i104,i106,i108,i110,i112,i114,i116,i118,i120,
i122,i124,i126,i128,i130,i132,i134,i136,i138,i140,i142,i144,i146,i148,i150,
i152,i154,i156,i158,i160,i162,i164,i166,i168,i170,i172,i174,i176,i178,i180,
i182,i184,i186,i188,i190,i192,i194,i196,i198,i200,i202,i204,i206,i208,i210,
i212,i214,i216,i218,i220,i222,i224,i226,i228,i230,i232,i234,i236,i238,i240,
i242,i244;

output p0,p1,p2,p3,p4,p5,p6,p7,p8,p9,p10,p11,p12,p13,p14,
p15,p16,p17,p18,p19,p20,p21,p22,p23,p24,p25,p26,p27,p28,p29,
p30,p31,p32,p33,p34,p35,p36,p37,p38,p39,p40,p41,p42,p43,p44,
p45,p46,p47,p48,p49,p50,p51,p52,p53,p54,p55,p56,p57,p58,p59,
p60,p61,p62,p63,p64,p65,p66,p67,p68,p69,p70,p71,p72,p73,p74,
p75,p76,p77,p78,p79,p80,p81,p82,p83,p84,p85,p86,p87,p88,p89,
p90,p91,p92,p93,p94,p95,p96,p97,p98,p99,p100,p101,p102,p103,p104,
p105,p106,p107,p108,p109,p110,p111,p112,p113,p114,p115,p116,p117,p118,p119,
p120,p121,p122,p123,p124,p125,p126,p127,p128,p129,p130,p131,p132,p133,p134,
p135,p136,p137,p138,p139,p140,p141,p142,p143,p144,p145,p146,p147,p148,p149,
p150,p151,p152,p153,p154,p155,p156,p157,p158,p159,p160,p161,p162,p163,p164,
p165,p166,p167,p168,p169,p170,p171,p172,p173,p174,p175,p176,p177,p178,p179,
p180,p181,p182,p183,p184,p185,p186,p187,p188,p189,p190,p191,p192,p193,p194,
p195,p196,p197,p198,p199,p200,p201,p202,p203,p204,p205,p206,p207,p208,p209,
p210,p211,p212,p213,p214,p215,p216,p217,p218,p219,p220,p221,p222,p223,p224,
p225,p226,p227,p228,p229,p230,p231,p232,p233,p234,p235,p236,p237,p238,p239,
p240,p241,p242,p243,p244,p245,p246,p247,p248,p249,p250,p251,p252,p253,p254,
p255,p256,p257,p258,p259,p260,p261,p262,p263,p264,p265,p266,p267,p268,p269,
p270,p271,p272,p273,p274,p275,p276,p277,p278,p279,p280,p281,p282,p283,p284,
p285,p286,p287,p288,p289,p290,p291,p292,p293,p294,p295,p296,p297,p298,p299,
p300,p301,p302,p303,p304,p305,p306,p307,p308,p309,p310,p311,p312,p313,p314,
p315,p316,p317,p318,p319,p320,p321,p322,p323,p324,p325,p326,p327,p328,p329,
p330,p331,p332,p333,p334,p335,p336,p337,p338,p339,p340,p341,p342,p343,p344,
p345,p346,p347,p348,p349,p350,p351,p352,p353,p354,p355,p356,p357,p358,p359,
p360,p361,p362,p363,p364,p365,p366,p367,p368,p369,p370,p371,p372,p373,p374,
p375,p376,p377,p378,p379,p380,p381,p382,p383,p384,p385,p386,p387,p388,p389,
p390,p391,p392,p393,p394,p395,p396,p397,p398,p399,p400,p401,p402,p403,p404,
p405,p406,p407,p408,p409,p410,p411,p412,p413,p414,p415,p416,p417,p418,p419,
p420,p421,p422,p423,p424,p425,p426,p427,p428,p429,p430,p431,p432,p433,p434,
p435,p436,p437,p438,p439,p440,p441,p442,p443,p444,p445,p446,p447,p448,p449,
p450,p451,p452,p453,p454,p455,p456,p457,p458,p459,p460,p461,p462,p463,p464,
p465,p466,p467,p468,p469,p470,p471,p472,p473,p474,p475,p476,p477,p478,p479,
p480,p481,p482,p483,p484,p485,p486,p487,p488,p489,p490,p491,p492,p493,p494,
p495,p496,p497,p498,p499,p500,p501,p502,p503,p504,p505,p506,p507,p508,p509,
p510,p511,p512,p513,p514,p515,p516,p517,p518,p519,p520,p521,p522,p523,p524,
p525,p526,p527,p528,p529,p530,p531,p532,p533,p534,p535,p536,p537,p538,p539,
p540,p541,p542,p543,p544,p545,p546,p547,p548,p549,p550,p551,p552,p553,p554,
p555,p556,p557,p558,p559,p560,p561,p562,p563,p564,p565,p566,p567,p568,p569,
p570,p571,p572,p573,p574,p575,p576,p577,p578,p579,p580,p581,p582,p583,p584,
p585,p586,p587,p588,p589,p590,p591,p592,p593,p594,p595,p596,p597,p598,p599,
p600,p601,p602,p603,p604,p605,p606,p607,p608,p609,p610,p611,p612,p613,p614,
p615,p616,p617,p618,p619,p620,p621,p622,p623,p624,p625,p626,p627,p628,p629,
p630,p631,p632,p633,p634,p635,p636,p637,p638,p639,p640,p641,p642,p643,p644,
p645,p646,p647,p648,p649,p650,p651,p652,p653,p654,p655,p656,p657,p658,p659,
p660,p661,p662,p663,p664,p665,p666,p667,p668,p669,p670,p671,p672,p673,p674,
p675,p676,p677,p678,p679,p680,p681,p682,p683,p684,p685,p686,p687,p688,p689,
p690,p691,p692,p693,p694,p695,p696,p697,p698,p699,p700,p701,p702,p703,p704,
p705,p706,p707,p708,p709,p710,p711,p712,p713,p714,p715,p716,p717,p718,p719,
p720,p721,p722,p723,p724,p725,p726,p727,p728,p729,p730,p731,p732,p733,p734,
p735,p736,p737,p738,p739,p740,p741,p742,p743,p744,p745,p746,p747,p748,p749,
p750,p751,p752,p753,p754,p755,p756,p757,p758,p759,p760,p761,p762,p763,p764,
p765,p766,p767,p768,p769,p770,p771,p772,p773,p774,p775,p776,p777,p778,p779,
p780,p781,p782,p783,p784,p785,p786,p787,p788,p789,p790,p791,p792,p793,p794,
p795,p796,p797,p798,p799,p800,p801,p802,p803,p804,p805,p806,p807,p808,p809,
p810,p811,p812,p813,p814,p815,p816,p817,p818,p819,p820,p821,p822,p823,p824,
p825,p826,p827,p828,p829,p830,p831,p832,p833,p834,p835,p836,p837,p838,p839,
p840,p841,p842,p843,p844,p845,p846,p847,p848,p849,p850,p851,p852,p853,p854,
p855,p856,p857,p858,p859,p860,p861,p862,p863,p864,p865,p866,p867,p868,p869,
p870,p871,p872,p873,p874,p875,p876,p877,p878,p879,p880,p881,p882,p883,p884,
p885,p886,p887,p888,p889,p890,p891,p892,p893,p894,p895,p896,p897,p898,p899,
p900,p901,p902,p903,p904,p905,p906,p907,p908,p909,p910,p911,p912,p913,p914,
p915,p916,p917,p918,p919,p920,p921,p922,p923,p924,p925,p926,p927,p928,p929,
p930,p931,p932,p933,p934,p935,p936,p937,p938,p939,p940,p941,p942,p943,p944,
p945,p946,p947,p948,p949,p950,p951,p952,p953,p954,p955,p956,p957,p958,p959,
p960,p961,p962,p963,p964,p965,p966,p967,p968,p969,p970,p971,p972,p973,p974,
p975,p976,p977,p978,p979,p980,p981,p982,p983,p984,p985,p986,p987,p988,p989,
p990,p991,p992,p993,p994,p995,p996,p997,p998,p999,p1000,p1001,p1002,p1003,p1004,
p1005,p1006,p1007,p1008,p1009,p1010,p1011,p1012,p1013,p1014,p1015,p1016,p1017,p1018,p1019,
p1020,p1021,p1022,p1023,p1024,p1025,p1026,p1027,p1028,p1029,p1030,p1031,p1032,p1033,p1034,
p1035,p1036,p1037,p1038,p1039,p1040,p1041,p1042,p1043,p1044,p1045,p1046,p1047,p1048,p1049,
p1050,p1051,p1052,p1053,p1054,p1055,p1056,p1057,p1058,p1059,p1060,p1061,p1062,p1063,p1064,
p1065,p1066,p1067,p1068,p1069,p1070,p1071,p1072,p1073,p1074,p1075,p1076,p1077,p1078,p1079,
p1080,p1081,p1082,p1083,p1084,p1085,p1086,p1087,p1088,p1089,p1090,p1091,p1092,p1093,p1094,
p1095,p1096,p1097,p1098,p1099,p1100,p1101,p1102,p1103,p1104,p1105,p1106,p1107,p1108,p1109,
p1110,p1111,p1112,p1113,p1114,p1115,p1116,p1117,p1118,p1119,p1120,p1121,p1122,p1123,p1124,
p1125,p1126,p1127,p1128,p1129,p1130,p1131,p1132,p1133,p1134,p1135,p1136,p1137,p1138,p1139,
p1140,p1141,p1142,p1143,p1144,p1145,p1146,p1147,p1148,p1149;

wire na2642,a2694,na2694,na2622,a2582,na2576,na2570,na2564,na2558,na2616,na2610,na2698,na2632,na2604,c1,
a2546,a2704,a2710,a2712,a2774,a2778,na2780,na2816,a2838,a2842,na2846,na2850,na2856,na2862,na2868,
na2874,na2880,na2886,na2892,na2898,na2904,na2908,a2910,a2916,a3060,a3080,a3200,na3230,a3232,na3238,
na3244,na3250,na3256,na3262,na3268,na3274,na3280,a3288,na3294,a3360,a3382,a3394,na3396,a3398,a3402,
na3410,na3420,na1206,a3428,a1228,a1314,na3438,a1316,a3448,a3452,a3456,na3460,na3486,na3498,a1230,
a3510,na3518,a3538,a3546,a3556,na2666,a3560,a3562,na3566,a3568,na3606,a3608,a3612,na3634,a3664,
na3734,na3770,a3794,na3820,a3824,a3826,na3836,a3842,a3848,a3854,a3860,a3866,a3872,a3878,a3884,
a3890,a3896,a3900,a1384,a1418,a3902,a3930,na1472,na3936,a3982,na1496,na4108,na4128,na4134,na4140,
na4146,a4158,na4174,na4180,na4186,na4192,na4202,na4224,na4238,na4244,na4250,na4256,na4262,na4290,na4304,
na4310,na4316,na4322,a4330,na4348,na4356,a4390,na4404,na4418,a4432,na4438,a4442,a4446,a4450,a4454,
a4458,a4462,a4466,a4470,a4474,a4478,na4480,a4486,a4492,a4498,na4504,a4514,a4520,a4526,na4534,
na4548,na4556,na4564,na4574,na4580,na4586,na4592,na4602,na4608,na4614,na4622,na4630,na4636,na4648,na4654,
na4660,na4666,na4672,na4678,na4684,na4690,na4696,na4702,na4710,na4716,na4722,na4728,na4734,na4740,na4746,
na4752,na4758,na4764,na4770,na4778,na4784,na4790,na4796,na4802,na4808,na4814,na4820,na4826,na4832,na4838,
na4844,na4850,na4856,na4862,na4868,na4874,na4880,na4886,na4892,na4898,na4904,na4910,na4916,na4922,na4928,
na4934,na4940,na4946,na4952,na4958,na4964,na4970,na4976,na4982,na4988,na4994,na5000,na5006,na5012,na5018,
na5024,na5030,na5036,na5042,na5048,na5054,na5060,na5066,na5072,na5078,na5084,na5090,na5096,na5102,na5108,
na5114,na5120,na5126,na5132,na5138,na5144,na5150,na5156,na5162,na5168,na5174,na5180,na5186,na5192,na5198,
na5204,na5210,na5216,na5222,na5228,na5234,na5240,na5244,a5250,na5262,na5274,na5286,a5296,a5298,a5300,
na5308,a5310,a5312,na5316,na5320,a5322,a5326,na5330,a5332,a5340,a5346,a5352,a5362,na5414,a5424,
na5442,a5444,a5450,na5456,a5464,a5472,a5480,a5492,a5500,a5510,a5518,a5526,a5534,a5540,a5546,
a5552,a5558,a5564,a5570,a5578,a5584,a5590,a5596,a5602,a5608,a5614,a5622,a5628,a5634,a5640,
a5646,a5652,a5660,a5666,a5672,a5678,a5684,a5690,a5696,a5704,a5710,a5716,a5722,a5728,a5734,
a5740,a5748,a5754,a5760,a5766,a5772,a5778,a5784,a5792,a5798,a5804,a5810,a5816,a5822,a5828,
na5830,a5834,a5888,a5918,a5948,a5978,a6008,na6102,a6106,a6110,a6112,a6114,a6116,na6138,na6148,
a1008,a1010,a1012,a1014,a1016,a1018,a1020,a1022,a1024,a1026,a1028,a1030,a1032,a1034,a1036,
a1038,a1040,a1042,a1044,a1046,a1048,a1050,a1052,a1054,a1056,a1058,a1060,a1062,a1064,a1066,
a1068,a1070,a1072,a1074,a1076,a1078,a1080,a1082,a1084,a1086,a1088,a1090,a1092,a1094,a1096,
a1098,a1100,a1102,a1104,a1106,a1108,a1110,a1112,a1114,a1116,a1118,a1120,a1122,a1124,a1126,
a1128,a1130,a1132,a1134,a1136,a1138,a1140,a1142,a1144,a1146,a1148,a1150,a1152,a1154,a1156,
a1158,a1160,a1162,a1164,a1166,a1168,a1170,a1172,a1174,a1176,a1178,a1180,a1182,a1184,a1186,
a1188,a1190,a1192,a1194,a1196,a1198,a1200,a1202,a1204,a1206,a1208,a1210,a1212,a1214,a1216,
a1218,a1220,a1222,a1224,a1226,a1232,a1234,a1236,a1238,a1240,a1242,a1244,a1246,a1248,a1250,
a1252,a1254,a1256,a1258,a1260,a1262,a1264,a1266,a1268,a1270,a1272,a1274,a1276,a1278,a1280,
a1282,a1284,a1286,a1288,a1290,a1292,a1294,a1296,a1298,a1300,a1302,a1304,a1306,a1308,a1310,
a1312,a1318,a1320,a1322,a1324,a1326,a1328,a1330,a1332,a1334,a1336,a1338,a1340,a1342,a1344,
a1346,a1348,a1350,a1352,a1354,a1356,a1358,a1360,a1362,a1364,a1366,a1368,a1370,a1372,a1374,
a1376,a1378,a1380,a1382,a1386,a1388,a1390,a1392,a1394,a1396,a1398,a1400,a1402,a1404,a1406,
a1408,a1410,a1412,a1414,a1416,a1420,a1422,a1424,a1426,a1428,a1430,a1432,a1434,a1436,a1438,
a1440,a1442,a1444,a1446,a1448,a1450,a1452,a1454,a1456,a1458,a1460,a1462,a1464,a1466,a1468,
a1470,a1472,a1474,a1476,a1478,a1480,a1482,a1484,a1486,a1488,a1490,a1492,a1494,a1496,a1498,
a1500,a1502,a1504,a1506,a1508,a1510,a1512,a1514,a1516,a1518,a1520,a1522,a1524,a1526,a1528,
a1530,a1532,a1534,a1536,a1538,a1540,a1542,a1544,a1546,a1548,a1550,a1552,a1554,a1556,a1558,
a1560,a1562,a1564,a1566,a1568,a1570,a1572,a1574,a1576,a1578,a1580,a1582,a1584,a1586,a1588,
a1590,a1592,a1594,a1596,a1598,a1600,a1602,a1604,a1606,a1608,a1610,a1612,a1614,a1616,a1618,
a1620,a1622,a1624,a1626,a1628,a1630,a1632,a1634,a1636,a1638,a1640,a1642,a1644,a1646,a1648,
a1650,a1652,a1654,a1656,a1658,a1660,a1662,a1664,a1666,a1668,a1670,a1672,a1674,a1676,a1678,
a1680,a1682,a1684,a1686,a1688,a1690,a1692,a1694,a1696,a1698,a1700,a1702,a1704,a1706,a1708,
a1710,a1712,a1714,a1716,a1718,a1720,a1722,a1724,a1726,a1728,a1730,a1732,a1734,a1736,a1738,
a1740,a1742,a1744,a1746,a1748,a1750,a1752,a1754,a1756,a1758,a1760,a1762,a1764,a1766,a1768,
a1770,a1772,a1774,a1776,a1778,a1780,a1782,a1784,a1786,a1788,a1790,a1792,a1794,a1796,a1798,
a1800,a1802,a1804,a1806,a1808,a1810,a1812,a1814,a1816,a1818,a1820,a1822,a1824,a1826,a1828,
a1830,a1832,a1834,a1836,a1838,a1840,a1842,a1844,a1846,a1848,a1850,a1852,a1854,a1856,a1858,
a1860,a1862,a1864,a1866,a1868,a1870,a1872,a1874,a1876,a1878,a1880,a1882,a1884,a1886,a1888,
a1890,a1892,a1894,a1896,a1898,a1900,a1902,a1904,a1906,a1908,a1910,a1912,a1914,a1916,a1918,
a1920,a1922,a1924,a1926,a1928,a1930,a1932,a1934,a1936,a1938,a1940,a1942,a1944,a1946,a1948,
a1950,a1952,a1954,a1956,a1958,a1960,a1962,a1964,a1966,a1968,a1970,a1972,a1974,a1976,a1978,
a1980,a1982,a1984,a1986,a1988,a1990,a1992,a1994,a1996,a1998,a2000,a2002,a2004,a2006,a2008,
a2010,a2012,a2014,a2016,a2018,a2020,a2022,a2024,a2026,a2028,a2030,a2032,a2034,a2036,a2038,
a2040,a2042,a2044,a2046,a2048,a2050,a2052,a2054,a2056,a2058,a2060,a2062,a2064,a2066,a2068,
a2070,a2072,a2074,a2076,a2078,a2080,a2082,a2084,a2086,a2088,a2090,a2092,a2094,a2096,a2098,
a2100,a2102,a2104,a2106,a2108,a2110,a2112,a2114,a2116,a2118,a2120,a2122,a2124,a2126,a2128,
a2130,a2132,a2134,a2136,a2138,a2140,a2142,a2144,a2146,a2148,a2150,a2152,a2154,a2156,a2158,
a2160,a2162,a2164,a2166,a2168,a2170,a2172,a2174,a2176,a2178,a2180,a2182,a2184,a2186,a2188,
a2190,a2192,a2194,a2196,a2198,a2200,a2202,a2204,a2206,a2208,a2210,a2212,a2214,a2216,a2218,
a2220,a2222,a2224,a2226,a2228,a2230,a2232,a2234,a2236,a2238,a2240,a2242,a2244,a2246,a2248,
a2250,a2252,a2254,a2256,a2258,a2260,a2262,a2264,a2266,a2268,a2270,a2272,a2274,a2276,a2278,
a2280,a2282,a2284,a2286,a2288,a2290,a2292,a2294,a2296,a2298,a2300,a2302,a2304,a2306,a2308,
a2310,a2312,a2314,a2316,a2318,a2320,a2322,a2324,a2326,a2328,a2330,a2332,a2334,a2336,a2338,
a2340,a2342,a2344,a2346,a2348,a2350,a2352,a2354,a2356,a2358,a2360,a2362,a2364,a2366,a2368,
a2370,a2372,a2374,a2376,a2378,a2380,a2382,a2384,a2386,a2388,a2390,a2392,a2394,a2396,a2398,
a2400,a2402,a2404,a2406,a2408,a2410,a2412,a2414,a2416,a2418,a2420,a2422,a2424,a2426,a2428,
a2430,a2432,a2434,a2436,a2438,a2440,a2442,a2444,a2446,a2448,a2450,a2452,a2454,a2456,a2458,
a2460,a2462,a2464,a2466,a2468,a2470,a2472,a2474,a2476,a2478,a2480,a2482,a2484,a2486,a2488,
a2490,a2492,a2494,a2496,a2498,a2500,a2502,a2504,a2506,a2508,a2510,a2512,a2514,a2516,a2518,
a2520,a2522,a2524,a2526,a2528,a2530,a2532,a2534,a2536,a2538,a2540,a2542,a2544,a2548,a2550,
a2552,a2554,a2556,a2558,a2560,a2562,a2564,a2566,a2568,a2570,a2572,a2574,a2576,a2578,a2580,
a2584,a2586,a2588,a2590,a2592,a2594,a2596,a2598,a2600,a2602,a2604,a2606,a2608,a2610,a2612,
a2614,a2616,a2618,a2620,a2622,a2624,a2626,a2628,a2630,a2632,a2634,a2636,a2638,a2640,a2642,
a2644,a2646,a2648,a2650,a2652,a2654,a2656,a2658,a2660,a2662,a2664,a2666,a2668,a2670,a2672,
a2674,a2676,a2678,a2680,a2682,a2684,a2686,a2688,a2690,a2692,a2696,a2698,a2700,a2702,a2706,
a2708,a2714,a2716,a2718,a2720,a2722,a2724,a2726,a2728,a2730,a2732,a2734,a2736,a2738,a2740,
a2742,a2744,a2746,a2748,a2750,a2752,a2754,a2756,a2758,a2760,a2762,a2764,a2766,a2768,a2770,
a2772,a2776,a2780,a2782,a2784,a2786,a2788,a2790,a2792,a2794,a2796,a2798,a2800,a2802,a2804,
a2806,a2808,a2810,a2812,a2814,a2816,a2818,a2820,a2822,a2824,a2826,a2828,a2830,a2832,a2834,
a2836,a2840,a2844,a2846,a2848,a2850,a2852,a2854,a2856,a2858,a2860,a2862,a2864,a2866,a2868,
a2870,a2872,a2874,a2876,a2878,a2880,a2882,a2884,a2886,a2888,a2890,a2892,a2894,a2896,a2898,
a2900,a2902,a2904,a2906,a2908,a2912,a2914,a2918,a2920,a2922,a2924,a2926,a2928,a2930,a2932,
a2934,a2936,a2938,a2940,a2942,a2944,a2946,a2948,a2950,a2952,a2954,a2956,a2958,a2960,a2962,
a2964,a2966,a2968,a2970,a2972,a2974,a2976,a2978,a2980,a2982,a2984,a2986,a2988,a2990,a2992,
a2994,a2996,a2998,a3000,a3002,a3004,a3006,a3008,a3010,a3012,a3014,a3016,a3018,a3020,a3022,
a3024,a3026,a3028,a3030,a3032,a3034,a3036,a3038,a3040,a3042,a3044,a3046,a3048,a3050,a3052,
a3054,a3056,a3058,a3062,a3064,a3066,a3068,a3070,a3072,a3074,a3076,a3078,a3082,a3084,a3086,
a3088,a3090,a3092,a3094,a3096,a3098,a3100,a3102,a3104,a3106,a3108,a3110,a3112,a3114,a3116,
a3118,a3120,a3122,a3124,a3126,a3128,a3130,a3132,a3134,a3136,a3138,a3140,a3142,a3144,a3146,
a3148,a3150,a3152,a3154,a3156,a3158,a3160,a3162,a3164,a3166,a3168,a3170,a3172,a3174,a3176,
a3178,a3180,a3182,a3184,a3186,a3188,a3190,a3192,a3194,a3196,a3198,a3202,a3204,a3206,a3208,
a3210,a3212,a3214,a3216,a3218,a3220,a3222,a3224,a3226,a3228,a3230,a3234,a3236,a3238,a3240,
a3242,a3244,a3246,a3248,a3250,a3252,a3254,a3256,a3258,a3260,a3262,a3264,a3266,a3268,a3270,
a3272,a3274,a3276,a3278,a3280,a3282,a3284,a3286,a3290,a3292,a3294,a3296,a3298,a3300,a3302,
a3304,a3306,a3308,a3310,a3312,a3314,a3316,a3318,a3320,a3322,a3324,a3326,a3328,a3330,a3332,
a3334,a3336,a3338,a3340,a3342,a3344,a3346,a3348,a3350,a3352,a3354,a3356,a3358,a3362,a3364,
a3366,a3368,a3370,a3372,a3374,a3376,a3378,a3380,a3384,a3386,a3388,a3390,a3392,a3396,a3400,
a3404,a3406,a3408,a3410,a3412,a3414,a3416,a3418,a3420,a3422,a3424,a3426,a3430,a3432,a3434,
a3436,a3438,a3440,a3442,a3444,a3446,a3450,a3454,a3458,a3460,a3462,a3464,a3466,a3468,a3470,
a3472,a3474,a3476,a3478,a3480,a3482,a3484,a3486,a3488,a3490,a3492,a3494,a3496,a3498,a3500,
a3502,a3504,a3506,a3508,a3512,a3514,a3516,a3518,a3520,a3522,a3524,a3526,a3528,a3530,a3532,
a3534,a3536,a3540,a3542,a3544,a3548,a3550,a3552,a3554,a3558,a3564,a3566,a3570,a3572,a3574,
a3576,a3578,a3580,a3582,a3584,a3586,a3588,a3590,a3592,a3594,a3596,a3598,a3600,a3602,a3604,
a3606,a3610,a3614,a3616,a3618,a3620,a3622,a3624,a3626,a3628,a3630,a3632,a3634,a3636,a3638,
a3640,a3642,a3644,a3646,a3648,a3650,a3652,a3654,a3656,a3658,a3660,a3662,a3666,a3668,a3670,
a3672,a3674,a3676,a3678,a3680,a3682,a3684,a3686,a3688,a3690,a3692,a3694,a3696,a3698,a3700,
a3702,a3704,a3706,a3708,a3710,a3712,a3714,a3716,a3718,a3720,a3722,a3724,a3726,a3728,a3730,
a3732,a3734,a3736,a3738,a3740,a3742,a3744,a3746,a3748,a3750,a3752,a3754,a3756,a3758,a3760,
a3762,a3764,a3766,a3768,a3770,a3772,a3774,a3776,a3778,a3780,a3782,a3784,a3786,a3788,a3790,
a3792,a3796,a3798,a3800,a3802,a3804,a3806,a3808,a3810,a3812,a3814,a3816,a3818,a3820,a3822,
a3828,a3830,a3832,a3834,a3836,a3838,a3840,a3844,a3846,a3850,a3852,a3856,a3858,a3862,a3864,
a3868,a3870,a3874,a3876,a3880,a3882,a3886,a3888,a3892,a3894,a3898,a3904,a3906,a3908,a3910,
a3912,a3914,a3916,a3918,a3920,a3922,a3924,a3926,a3928,a3932,a3934,a3936,a3938,a3940,a3942,
a3944,a3946,a3948,a3950,a3952,a3954,a3956,a3958,a3960,a3962,a3964,a3966,a3968,a3970,a3972,
a3974,a3976,a3978,a3980,a3984,a3986,a3988,a3990,a3992,a3994,a3996,a3998,a4000,a4002,a4004,
a4006,a4008,a4010,a4012,a4014,a4016,a4018,a4020,a4022,a4024,a4026,a4028,a4030,a4032,a4034,
a4036,a4038,a4040,a4042,a4044,a4046,a4048,a4050,a4052,a4054,a4056,a4058,a4060,a4062,a4064,
a4066,a4068,a4070,a4072,a4074,a4076,a4078,a4080,a4082,a4084,a4086,a4088,a4090,a4092,a4094,
a4096,a4098,a4100,a4102,a4104,a4106,a4108,a4110,a4112,a4114,a4116,a4118,a4120,a4122,a4124,
a4126,a4128,a4130,a4132,a4134,a4136,a4138,a4140,a4142,a4144,a4146,a4148,a4150,a4152,a4154,
a4156,a4160,a4162,a4164,a4166,a4168,a4170,a4172,a4174,a4176,a4178,a4180,a4182,a4184,a4186,
a4188,a4190,a4192,a4194,a4196,a4198,a4200,a4202,a4204,a4206,a4208,a4210,a4212,a4214,a4216,
a4218,a4220,a4222,a4224,a4226,a4228,a4230,a4232,a4234,a4236,a4238,a4240,a4242,a4244,a4246,
a4248,a4250,a4252,a4254,a4256,a4258,a4260,a4262,a4264,a4266,a4268,a4270,a4272,a4274,a4276,
a4278,a4280,a4282,a4284,a4286,a4288,a4290,a4292,a4294,a4296,a4298,a4300,a4302,a4304,a4306,
a4308,a4310,a4312,a4314,a4316,a4318,a4320,a4322,a4324,a4326,a4328,a4332,a4334,a4336,a4338,
a4340,a4342,a4344,a4346,a4348,a4350,a4352,a4354,a4356,a4358,a4360,a4362,a4364,a4366,a4368,
a4370,a4372,a4374,a4376,a4378,a4380,a4382,a4384,a4386,a4388,a4392,a4394,a4396,a4398,a4400,
a4402,a4404,a4406,a4408,a4410,a4412,a4414,a4416,a4418,a4420,a4422,a4424,a4426,a4428,a4430,
a4434,a4436,a4438,a4440,a4444,a4448,a4452,a4456,a4460,a4464,a4468,a4472,a4476,a4480,a4482,
a4484,a4488,a4490,a4494,a4496,a4500,a4502,a4504,a4506,a4508,a4510,a4512,a4516,a4518,a4522,
a4524,a4528,a4530,a4532,a4534,a4536,a4538,a4540,a4542,a4544,a4546,a4548,a4550,a4552,a4554,
a4556,a4558,a4560,a4562,a4564,a4566,a4568,a4570,a4572,a4574,a4576,a4578,a4580,a4582,a4584,
a4586,a4588,a4590,a4592,a4594,a4596,a4598,a4600,a4602,a4604,a4606,a4608,a4610,a4612,a4614,
a4616,a4618,a4620,a4622,a4624,a4626,a4628,a4630,a4632,a4634,a4636,a4638,a4640,a4642,a4644,
a4646,a4648,a4650,a4652,a4654,a4656,a4658,a4660,a4662,a4664,a4666,a4668,a4670,a4672,a4674,
a4676,a4678,a4680,a4682,a4684,a4686,a4688,a4690,a4692,a4694,a4696,a4698,a4700,a4702,a4704,
a4706,a4708,a4710,a4712,a4714,a4716,a4718,a4720,a4722,a4724,a4726,a4728,a4730,a4732,a4734,
a4736,a4738,a4740,a4742,a4744,a4746,a4748,a4750,a4752,a4754,a4756,a4758,a4760,a4762,a4764,
a4766,a4768,a4770,a4772,a4774,a4776,a4778,a4780,a4782,a4784,a4786,a4788,a4790,a4792,a4794,
a4796,a4798,a4800,a4802,a4804,a4806,a4808,a4810,a4812,a4814,a4816,a4818,a4820,a4822,a4824,
a4826,a4828,a4830,a4832,a4834,a4836,a4838,a4840,a4842,a4844,a4846,a4848,a4850,a4852,a4854,
a4856,a4858,a4860,a4862,a4864,a4866,a4868,a4870,a4872,a4874,a4876,a4878,a4880,a4882,a4884,
a4886,a4888,a4890,a4892,a4894,a4896,a4898,a4900,a4902,a4904,a4906,a4908,a4910,a4912,a4914,
a4916,a4918,a4920,a4922,a4924,a4926,a4928,a4930,a4932,a4934,a4936,a4938,a4940,a4942,a4944,
a4946,a4948,a4950,a4952,a4954,a4956,a4958,a4960,a4962,a4964,a4966,a4968,a4970,a4972,a4974,
a4976,a4978,a4980,a4982,a4984,a4986,a4988,a4990,a4992,a4994,a4996,a4998,a5000,a5002,a5004,
a5006,a5008,a5010,a5012,a5014,a5016,a5018,a5020,a5022,a5024,a5026,a5028,a5030,a5032,a5034,
a5036,a5038,a5040,a5042,a5044,a5046,a5048,a5050,a5052,a5054,a5056,a5058,a5060,a5062,a5064,
a5066,a5068,a5070,a5072,a5074,a5076,a5078,a5080,a5082,a5084,a5086,a5088,a5090,a5092,a5094,
a5096,a5098,a5100,a5102,a5104,a5106,a5108,a5110,a5112,a5114,a5116,a5118,a5120,a5122,a5124,
a5126,a5128,a5130,a5132,a5134,a5136,a5138,a5140,a5142,a5144,a5146,a5148,a5150,a5152,a5154,
a5156,a5158,a5160,a5162,a5164,a5166,a5168,a5170,a5172,a5174,a5176,a5178,a5180,a5182,a5184,
a5186,a5188,a5190,a5192,a5194,a5196,a5198,a5200,a5202,a5204,a5206,a5208,a5210,a5212,a5214,
a5216,a5218,a5220,a5222,a5224,a5226,a5228,a5230,a5232,a5234,a5236,a5238,a5240,a5242,a5244,
a5246,a5248,a5252,a5254,a5256,a5258,a5260,a5262,a5264,a5266,a5268,a5270,a5272,a5274,a5276,
a5278,a5280,a5282,a5284,a5286,a5288,a5290,a5292,a5294,a5302,a5304,a5306,a5308,a5314,a5316,
a5318,a5320,a5324,a5328,a5330,a5334,a5336,a5338,a5342,a5344,a5348,a5350,a5354,a5356,a5358,
a5360,a5364,a5366,a5368,a5370,a5372,a5374,a5376,a5378,a5380,a5382,a5384,a5386,a5388,a5390,
a5392,a5394,a5396,a5398,a5400,a5402,a5404,a5406,a5408,a5410,a5412,a5414,a5416,a5418,a5420,
a5422,a5426,a5428,a5430,a5432,a5434,a5436,a5438,a5440,a5442,a5446,a5448,a5452,a5454,a5456,
a5458,a5460,a5462,a5466,a5468,a5470,a5474,a5476,a5478,a5482,a5484,a5486,a5488,a5490,a5494,
a5496,a5498,a5502,a5504,a5506,a5508,a5512,a5514,a5516,a5520,a5522,a5524,a5528,a5530,a5532,
a5536,a5538,a5542,a5544,a5548,a5550,a5554,a5556,a5560,a5562,a5566,a5568,a5572,a5574,a5576,
a5580,a5582,a5586,a5588,a5592,a5594,a5598,a5600,a5604,a5606,a5610,a5612,a5616,a5618,a5620,
a5624,a5626,a5630,a5632,a5636,a5638,a5642,a5644,a5648,a5650,a5654,a5656,a5658,a5662,a5664,
a5668,a5670,a5674,a5676,a5680,a5682,a5686,a5688,a5692,a5694,a5698,a5700,a5702,a5706,a5708,
a5712,a5714,a5718,a5720,a5724,a5726,a5730,a5732,a5736,a5738,a5742,a5744,a5746,a5750,a5752,
a5756,a5758,a5762,a5764,a5768,a5770,a5774,a5776,a5780,a5782,a5786,a5788,a5790,a5794,a5796,
a5800,a5802,a5806,a5808,a5812,a5814,a5818,a5820,a5824,a5826,a5830,a5832,a5836,a5838,a5840,
a5842,a5844,a5846,a5848,a5850,a5852,a5854,a5856,a5858,a5860,a5862,a5864,a5866,a5868,a5870,
a5872,a5874,a5876,a5878,a5880,a5882,a5884,a5886,a5890,a5892,a5894,a5896,a5898,a5900,a5902,
a5904,a5906,a5908,a5910,a5912,a5914,a5916,a5920,a5922,a5924,a5926,a5928,a5930,a5932,a5934,
a5936,a5938,a5940,a5942,a5944,a5946,a5950,a5952,a5954,a5956,a5958,a5960,a5962,a5964,a5966,
a5968,a5970,a5972,a5974,a5976,a5980,a5982,a5984,a5986,a5988,a5990,a5992,a5994,a5996,a5998,
a6000,a6002,a6004,a6006,a6010,a6012,a6014,a6016,a6018,a6020,a6022,a6024,a6026,a6028,a6030,
a6032,a6034,a6036,a6038,a6040,a6042,a6044,a6046,a6048,a6050,a6052,a6054,a6056,a6058,a6060,
a6062,a6064,a6066,a6068,a6070,a6072,a6074,a6076,a6078,a6080,a6082,a6084,a6086,a6088,a6090,
a6092,a6094,a6096,a6098,a6100,a6102,a6104,a6108,a6118,a6120,a6122,a6124,a6126,a6128,a6130,
a6132,a6134,a6136,a6138,a6140,a6142,a6144,a6146,a6148,p0,c0,p1,p2,p3,p4,
p5,p6,p7,p8,p9,p10,p11,p12,p13,p14,p15,p16,p17,p18,p19,
p20,p21,p22,p23,p24,p25,p26,p27,p28,p29,p30,p31,p32,p33,p34,
p35,p36,p37,p38,p39,p40,p41,p42,p43,p44,p45,p46,p47,p48,p49,
p50,p51,p52,p53,p54,p55,p56,p57,p58,p59,p60,p61,p62,p63,p64,
p65,p66,p67,p68,p69,p70,p71,p72,p73,p74,p75,p76,p77,p78,p79,
p80,p81,p82,p83,p84,p85,p86,p87,p88,p89,p90,p91,p92,p93,p94,
p95,p96,p97,p98,p99,p100,p101,p102,p103,p104,p105,p106,p107,p108,p109,
p110,p111,p112,p113,p114,p115,p116,p117,p118,p119,p120,p121,p122,p123,p124,
p125,p126,p127,p128,p129,p130,p131,p132,p133,p134,p135,p136,p137,p138,p139,
p140,p141,p142,p143,p144,p145,p146,p147,p148,p149,p150,p151,p152,p153,p154,
p155,p156,p157,p158,p159,p160,p161,p162,p163,p164,p165,p166,p167,p168,p169,
p170,p171,p172,p173,p174,p175,p176,p177,p178,p179,p180,p181,p182,p183,p184,
p185,p186,p187,p188,p189,p190,p191,p192,p193,p194,p195,p196,p197,p198,p199,
p200,p201,p202,p203,p204,p205,p206,p207,p208,p209,p210,p211,p212,p213,p214,
p215,p216,p217,p218,p219,p220,p221,p222,p223,p224,p225,p226,p227,p228,p229,
p230,p231,p232,p233,p234,p235,p236,p237,p238,p239,p240,p241,p242,p243,p244,
p245,p246,p247,p248,p249,p250,p251,p252,p253,p254,p255,p256,p257,p258,p259,
p260,p261,p262,p263,p264,p265,p266,p267,p268,p269,p270,p271,p272,p273,p274,
p275,p276,p277,p278,p279,p280,p281,p282,p283,p284,p285,p286,p287,p288,p289,
p290,p291,p292,p293,p294,p295,p296,p297,p298,p299,p300,p301,p302,p303,p304,
p305,p306,p307,p308,p309,p310,p311,p312,p313,p314,p315,p316,p317,p318,p319,
p320,p321,p322,p323,p324,p325,p326,p327,p328,p329,p330,p331,p332,p333,p334,
p335,p336,p337,p338,p339,p340,p341,p342,p343,p344,p345,p346,p347,p348,p349,
p350,p351,p352,p353,p354,p355,p356,p357,p358,p359,p360,p361,p362,p363,p364,
p365,p366,p367,p368,p369,p370,p371,p372,p373,p374,p375,p376,p377,p378,p379,
p380,p381,p382,p383,p384,p385,p386,p387,p388,p389,p390,p391,p392,p393,p394,
p395,p396,p397,p398,p399,p400,p401,p402,p403,p404,p405,p406,p407,p408,p409,
p410,p411,p412,p413,p414,p415,p416,p417,p418,p419,p420,p421,p422,p423,p424,
p425,p426,p427,p428,p429,p430,p431,p432,p433,p434,p435,p436,p437,p438,p439,
p440,p441,p442,p443,p444,p445,p446,p447,p448,p449,p450,p451,p452,p453,p454,
p455,p456,p457,p458,p459,p460,p461,p462,p463,p464,p465,p466,p467,p468,p469,
p470,p471,p472,p473,p474,p475,p476,p477,p478,p479,p480,p481,p482,p483,p484,
p485,p486,p487,p488,p489,p490,p491,p492,p493,p494,p495,p496,p497,p498,p499,
p500,p501,p502,p503,p504,p505,p506,p507,p508,p509,p510,p511,p512,p513,p514,
p515,p516,p517,p518,p519,p520,p521,p522,p523,p524,p525,p526,p527,p528,p529,
p530,p531,p532,p533,p534,p535,p536,p537,p538,p539,p540,p541,p542,p543,p544,
p545,p546,p547,p548,p549,p550,p551,p552,p553,p554,p555,p556,p557,p558,p559,
p560,p561,p562,p563,p564,p565,p566,p567,p568,p569,p570,p571,p572,p573,p574,
p575,p576,p577,p578,p579,p580,p581,p582,p583,p584,p585,p586,p587,p588,p589,
p590,p591,p592,p593,p594,p595,p596,p597,p598,p599,p600,p601,p602,p603,p604,
p605,p606,p607,p608,p609,p610,p611,p612,p613,p614,p615,p616,p617,p618,p619,
p620,p621,p622,p623,p624,p625,p626,p627,p628,p629,p630,p631,p632,p633,p634,
p635,p636,p637,p638,p639,p640,p641,p642,p643,p644,p645,p646,p647,p648,p649,
p650,p651,p652,p653,p654,p655,p656,p657,p658,p659,p660,p661,p662,p663,p664,
p665,p666,p667,p668,p669,p670,p671,p672,p673,p674,p675,p676,p677,p678,p679,
p680,p681,p682,p683,p684,p685,p686,p687,p688,p689,p690,p691,p692,p693,p694,
p695,p696,p697,p698,p699,p700,p701,p702,p703,p704,p705,p706,p707,p708,p709,
p710,p711,p712,p713,p714,p715,p716,p717,p718,p719,p720,p721,p722,p723,p724,
p725,p726,p727,p728,p729,p730,p731,p732,p733,p734,p735,p736,p737,p738,p739,
p740,p741,p742,p743,p744,p745,p746,p747,p748,p749,p750,p751,p752,p753,p754,
p755,p756,p757,p758,p759,p760,p761,p762,p763,p764,p765,p766,p767,p768,p769,
p770,p771,p772,p773,p774,p775,p776,p777,p778,p779,p780,p781,p782,p783,p784,
p785,p786,p787,p788,p789,p790,p791,p792,p793,p794,p795,p796,p797,p798,p799,
p800,p801,p802,p803,p804,p805,p806,p807,p808,p809,p810,p811,p812,p813,p814,
p815,p816,p817,p818,p819,p820,p821,p822,p823,p824,p825,p826,p827,p828,p829,
p830,p831,p832,p833,p834,p835,p836,p837,p838,p839,p840,p841,p842,p843,p844,
p845,p846,p847,p848,p849,p850,p851,p852,p853,p854,p855,p856,p857,p858,p859,
p860,p861,p862,p863,p864,p865,p866,p867,p868,p869,p870,p871,p872,p873,p874,
p875,p876,p877,p878,p879,p880,p881,p882,p883,p884,p885,p886,p887,p888,p889,
p890,p891,p892,p893,p894,p895,p896,p897,p898,p899,p900,p901,p902,p903,p904,
p905,p906,p907,p908,p909,p910,p911,p912,p913,p914,p915,p916,p917,p918,p919,
p920,p921,p922,p923,p924,p925,p926,p927,p928,p929,p930,p931,p932,p933,p934,
p935,p936,p937,p938,p939,p940,p941,p942,p943,p944,p945,p946,p947,p948,p949,
p950,p951,p952,p953,p954,p955,p956,p957,p958,p959,p960,p961,p962,p963,p964,
p965,p966,p967,p968,p969,p970,p971,p972,p973,p974,p975,p976,p977,p978,p979,
p980,p981,p982,p983,p984,p985,p986,p987,p988,p989,p990,p991,p992,p993,p994,
p995,p996,p997,p998,p999,p1000,p1001,p1002,p1003,p1004,p1005,p1006,p1007,p1008,p1009,
p1010,p1011,p1012,p1013,p1014,p1015,p1016,p1017,p1018,p1019,p1020,p1021,p1022,p1023,p1024,
p1025,p1026,p1027,p1028,p1029,p1030,p1031,p1032,p1033,p1034,p1035,p1036,p1037,p1038,p1039,
p1040,p1041,p1042,p1043,p1044,p1045,p1046,p1047,p1048,p1049,p1050,p1051,p1052,p1053,p1054,
p1055,p1056,p1057,p1058,p1059,p1060,p1061,p1062,p1063,p1064,p1065,p1066,p1067,p1068,p1069,
p1070,p1071,p1072,p1073,p1074,p1075,p1076,p1077,p1078,p1079,p1080,p1081,p1082,p1083,p1084,
p1085,p1086,p1087,p1088,p1089,p1090,p1091,p1092,p1093,p1094,p1095,p1096,p1097,p1098,p1099,
p1100,p1101,p1102,p1103,p1104,p1105,p1106,p1107,p1108,p1109,p1110,p1111,p1112,p1113,p1114,
p1115,p1116,p1117,p1118,p1119,p1120,p1121,p1122,p1123,p1124,p1125,p1126,p1127,p1128,p1129,
p1130,p1131,p1132,p1133,p1134,p1135,p1136,p1137,p1138,p1139,p1140,p1141,p1142,p1143,p1144,
p1145,p1146,p1147,p1148,p1149;

reg l246,l248,l250,l252,l254,l256,l258,l260,l262,l264,l266,l268,l270,l272,l274,
l276,l278,l280,l282,l284,l286,l288,l290,l292,l294,l296,l298,l300,l302,l304,
l306,l308,l310,l312,l314,l316,l318,l320,l322,l324,l326,l328,l330,l332,l334,
l336,l338,l340,l342,l344,l346,l348,l350,l352,l354,l356,l358,l360,l362,l364,
l366,l368,l370,l372,l374,l376,l378,l380,l382,l384,l386,l388,l390,l392,l394,
l396,l398,l400,l402,l404,l406,l408,l410,l412,l414,l416,l418,l420,l422,l424,
l426,l428,l430,l432,l434,l436,l438,l440,l442,l444,l446,l448,l450,l452,l454,
l456,l458,l460,l462,l464,l466,l468,l470,l472,l474,l476,l478,l480,l482,l484,
l486,l488,l490,l492,l494,l496,l498,l500,l502,l504,l506,l508,l510,l512,l514,
l516,l518,l520,l522,l524,l526,l528,l530,l532,l534,l536,l538,l540,l542,l544,
l546,l548,l550,l552,l554,l556,l558,l560,l562,l564,l566,l568,l570,l572,l574,
l576,l578,l580,l582,l584,l586,l588,l590,l592,l594,l596,l598,l600,l602,l604,
l606,l608,l610,l612,l614,l616,l618,l620,l622,l624,l626,l628,l630,l632,l634,
l636,l638,l640,l642,l644,l646,l648,l650,l652,l654,l656,l658,l660,l662,l664,
l666,l668,l670,l672,l674,l676,l678,l680,l682,l684,l686,l688,l690,l692,l694,
l696,l698,l700,l702,l704,l706,l708,l710,l712,l714,l716,l718,l720,l722,l724,
l726,l728,l730,l732,l734,l736,l738,l740,l742,l744,l746,l748,l750,l752,l754,
l756,l758,l760,l762,l764,l766,l768,l770,l772,l774,l776,l778,l780,l782,l784,
l786,l788,l790,l792,l794,l796,l798,l800,l802,l804,l806,l808,l810,l812,l814,
l816,l818,l820,l822,l824,l826,l828,l830,l832,l834,l836,l838,l840,l842,l844,
l846,l848,l850,l852,l854,l856,l858,l860,l862,l864,l866,l868,l870,l872,l874,
l876,l878,l880,l882,l884,l886,l888,l890,l892,l894,l896,l898,l900,l902,l904,
l906,l908,l910,l912,l914,l916,l918,l920,l922,l924,l926,l928,l930,l932,l934,
l936,l938,l940,l942,l944,l946,l948,l950,l952,l954,l956,l958,l960,l962,l964,
l966,l968,l970,l972,l974,l976,l978,l980,l982,l984,l986,l988,l990,l992,l994,
l996,l998,l1000,l1002,l1004,l1006;

initial
begin
   l246 = 0;
   l248 = 0;
   l250 = 0;
   l252 = 0;
   l254 = 0;
   l256 = 0;
   l258 = 0;
   l260 = 0;
   l262 = 0;
   l264 = 0;
   l266 = 0;
   l268 = 0;
   l270 = 0;
   l272 = 0;
   l274 = 0;
   l276 = 0;
   l278 = 0;
   l280 = 0;
   l282 = 0;
   l284 = 0;
   l286 = 0;
   l288 = 0;
   l290 = 0;
   l292 = 0;
   l294 = 0;
   l296 = 0;
   l298 = 0;
   l300 = 0;
   l302 = 0;
   l304 = 0;
   l306 = 0;
   l308 = 0;
   l310 = 0;
   l312 = 0;
   l314 = 0;
   l316 = 0;
   l318 = 0;
   l320 = 0;
   l322 = 0;
   l324 = 0;
   l326 = 0;
   l328 = 0;
   l330 = 0;
   l332 = 0;
   l334 = 0;
   l336 = 0;
   l338 = 0;
   l340 = 0;
   l342 = 0;
   l344 = 0;
   l346 = 0;
   l348 = 0;
   l350 = 0;
   l352 = 0;
   l354 = 0;
   l356 = 0;
   l358 = 0;
   l360 = 0;
   l362 = 0;
   l364 = 0;
   l366 = 0;
   l368 = 0;
   l370 = 0;
   l372 = 0;
   l374 = 0;
   l376 = 0;
   l378 = 0;
   l380 = 0;
   l382 = 0;
   l384 = 0;
   l386 = 0;
   l388 = 0;
   l390 = 0;
   l392 = 0;
   l394 = 0;
   l396 = 0;
   l398 = 0;
   l400 = 0;
   l402 = 0;
   l404 = 0;
   l406 = 0;
   l408 = 0;
   l410 = 0;
   l412 = 0;
   l414 = 0;
   l416 = 0;
   l418 = 0;
   l420 = 0;
   l422 = 0;
   l424 = 0;
   l426 = 0;
   l428 = 0;
   l430 = 0;
   l432 = 0;
   l434 = 0;
   l436 = 0;
   l438 = 0;
   l440 = 0;
   l442 = 0;
   l444 = 0;
   l446 = 0;
   l448 = 0;
   l450 = 0;
   l452 = 0;
   l454 = 0;
   l456 = 0;
   l458 = 0;
   l460 = 0;
   l462 = 0;
   l464 = 0;
   l466 = 0;
   l468 = 0;
   l470 = 0;
   l472 = 0;
   l474 = 0;
   l476 = 0;
   l478 = 0;
   l480 = 0;
   l482 = 0;
   l484 = 0;
   l486 = 0;
   l488 = 0;
   l490 = 0;
   l492 = 0;
   l494 = 0;
   l496 = 0;
   l498 = 0;
   l500 = 0;
   l502 = 0;
   l504 = 0;
   l506 = 0;
   l508 = 0;
   l510 = 0;
   l512 = 0;
   l514 = 0;
   l516 = 0;
   l518 = 0;
   l520 = 0;
   l522 = 0;
   l524 = 0;
   l526 = 0;
   l528 = 0;
   l530 = 0;
   l532 = 0;
   l534 = 0;
   l536 = 0;
   l538 = 0;
   l540 = 0;
   l542 = 0;
   l544 = 0;
   l546 = 0;
   l548 = 0;
   l550 = 0;
   l552 = 0;
   l554 = 0;
   l556 = 0;
   l558 = 0;
   l560 = 0;
   l562 = 0;
   l564 = 0;
   l566 = 0;
   l568 = 0;
   l570 = 0;
   l572 = 0;
   l574 = 0;
   l576 = 0;
   l578 = 0;
   l580 = 0;
   l582 = 0;
   l584 = 0;
   l586 = 0;
   l588 = 0;
   l590 = 0;
   l592 = 0;
   l594 = 0;
   l596 = 0;
   l598 = 0;
   l600 = 0;
   l602 = 0;
   l604 = 0;
   l606 = 0;
   l608 = 0;
   l610 = 0;
   l612 = 0;
   l614 = 0;
   l616 = 0;
   l618 = 0;
   l620 = 0;
   l622 = 0;
   l624 = 0;
   l626 = 0;
   l628 = 0;
   l630 = 0;
   l632 = 0;
   l634 = 0;
   l636 = 0;
   l638 = 0;
   l640 = 0;
   l642 = 0;
   l644 = 0;
   l646 = 0;
   l648 = 0;
   l650 = 0;
   l652 = 0;
   l654 = 0;
   l656 = 0;
   l658 = 0;
   l660 = 0;
   l662 = 0;
   l664 = 0;
   l666 = 0;
   l668 = 0;
   l670 = 0;
   l672 = 0;
   l674 = 0;
   l676 = 0;
   l678 = 0;
   l680 = 0;
   l682 = 0;
   l684 = 0;
   l686 = 0;
   l688 = 0;
   l690 = 0;
   l692 = 0;
   l694 = 0;
   l696 = 0;
   l698 = 0;
   l700 = 0;
   l702 = 0;
   l704 = 0;
   l706 = 0;
   l708 = 0;
   l710 = 0;
   l712 = 0;
   l714 = 0;
   l716 = 0;
   l718 = 0;
   l720 = 0;
   l722 = 0;
   l724 = 0;
   l726 = 0;
   l728 = 0;
   l730 = 0;
   l732 = 0;
   l734 = 0;
   l736 = 0;
   l738 = 0;
   l740 = 0;
   l742 = 0;
   l744 = 0;
   l746 = 0;
   l748 = 0;
   l750 = 0;
   l752 = 0;
   l754 = 0;
   l756 = 0;
   l758 = 0;
   l760 = 0;
   l762 = 0;
   l764 = 0;
   l766 = 0;
   l768 = 0;
   l770 = 0;
   l772 = 0;
   l774 = 0;
   l776 = 0;
   l778 = 0;
   l780 = 0;
   l782 = 0;
   l784 = 0;
   l786 = 0;
   l788 = 0;
   l790 = 0;
   l792 = 0;
   l794 = 0;
   l796 = 0;
   l798 = 0;
   l800 = 0;
   l802 = 0;
   l804 = 0;
   l806 = 0;
   l808 = 0;
   l810 = 0;
   l812 = 0;
   l814 = 0;
   l816 = 0;
   l818 = 0;
   l820 = 0;
   l822 = 0;
   l824 = 0;
   l826 = 0;
   l828 = 0;
   l830 = 0;
   l832 = 0;
   l834 = 0;
   l836 = 0;
   l838 = 0;
   l840 = 0;
   l842 = 0;
   l844 = 0;
   l846 = 0;
   l848 = 0;
   l850 = 0;
   l852 = 0;
   l854 = 0;
   l856 = 0;
   l858 = 0;
   l860 = 0;
   l862 = 0;
   l864 = 0;
   l866 = 0;
   l868 = 0;
   l870 = 0;
   l872 = 0;
   l874 = 0;
   l876 = 0;
   l878 = 0;
   l880 = 0;
   l882 = 0;
   l884 = 0;
   l886 = 0;
   l888 = 0;
   l890 = 0;
   l892 = 0;
   l894 = 0;
   l896 = 0;
   l898 = 0;
   l900 = 0;
   l902 = 0;
   l904 = 0;
   l906 = 0;
   l908 = 0;
   l910 = 0;
   l912 = 0;
   l914 = 0;
   l916 = 0;
   l918 = 0;
   l920 = 0;
   l922 = 0;
   l924 = 0;
   l926 = 0;
   l928 = 0;
   l930 = 0;
   l932 = 0;
   l934 = 0;
   l936 = 0;
   l938 = 0;
   l940 = 0;
   l942 = 0;
   l944 = 0;
   l946 = 0;
   l948 = 0;
   l950 = 0;
   l952 = 0;
   l954 = 0;
   l956 = 0;
   l958 = 0;
   l960 = 0;
   l962 = 0;
   l964 = 0;
   l966 = 0;
   l968 = 0;
   l970 = 0;
   l972 = 0;
   l974 = 0;
   l976 = 0;
   l978 = 0;
   l980 = 0;
   l982 = 0;
   l984 = 0;
   l986 = 0;
   l988 = 0;
   l990 = 0;
   l992 = 0;
   l994 = 0;
   l996 = 0;
   l998 = 0;
   l1000 = 0;
   l1002 = 0;
   l1004 = 0;
   l1006 = 0;
end

always @(posedge na2642)
   l246 <= na2642;

always @(posedge a2694)
   l248 <= a2694;

always @(posedge na2694)
   l250 <= na2694;

always @(posedge na2622)
   l252 <= na2622;

always @(posedge a2582)
   l254 <= a2582;

always @(posedge na2576)
   l256 <= na2576;

always @(posedge na2570)
   l258 <= na2570;

always @(posedge na2564)
   l260 <= na2564;

always @(posedge na2558)
   l262 <= na2558;

always @(posedge na2616)
   l264 <= na2616;

always @(posedge na2610)
   l266 <= na2610;

always @(posedge na2698)
   l268 <= na2698;

always @(posedge na2632)
   l270 <= na2632;

always @(posedge na2604)
   l272 <= na2604;

always @(posedge c1)
   l274 <= c1;

always @(posedge l370)
   l276 <= l370;

always @(posedge l420)
   l278 <= l420;

always @(posedge l858)
   l280 <= l858;

always @(posedge l982)
   l282 <= l982;

always @(posedge a2546)
   l284 <= a2546;

always @(posedge l1000)
   l286 <= l1000;

always @(posedge a2704)
   l288 <= a2704;

always @(posedge a2710)
   l290 <= a2710;

always @(posedge a2712)
   l292 <= a2712;

always @(posedge a2774)
   l294 <= a2774;

always @(posedge a2778)
   l296 <= a2778;

always @(posedge na2780)
   l298 <= na2780;

always @(posedge na2816)
   l300 <= na2816;

always @(posedge a2838)
   l302 <= a2838;

always @(posedge a2842)
   l304 <= a2842;

always @(posedge na2846)
   l306 <= na2846;

always @(posedge na2850)
   l308 <= na2850;

always @(posedge na2856)
   l310 <= na2856;

always @(posedge na2862)
   l312 <= na2862;

always @(posedge na2868)
   l314 <= na2868;

always @(posedge na2874)
   l316 <= na2874;

always @(posedge na2880)
   l318 <= na2880;

always @(posedge na2886)
   l320 <= na2886;

always @(posedge na2892)
   l322 <= na2892;

always @(posedge na2898)
   l324 <= na2898;

always @(posedge na2904)
   l326 <= na2904;

always @(posedge na2908)
   l328 <= na2908;

always @(posedge a2910)
   l330 <= a2910;

always @(posedge a2916)
   l332 <= a2916;

always @(posedge a3060)
   l334 <= a3060;

always @(posedge a3080)
   l336 <= a3080;

always @(posedge a3200)
   l338 <= a3200;

always @(posedge na3230)
   l340 <= na3230;

always @(posedge a3232)
   l342 <= a3232;

always @(posedge na3238)
   l344 <= na3238;

always @(posedge na3244)
   l346 <= na3244;

always @(posedge na3250)
   l348 <= na3250;

always @(posedge na3256)
   l350 <= na3256;

always @(posedge na3262)
   l352 <= na3262;

always @(posedge na3268)
   l354 <= na3268;

always @(posedge na3274)
   l356 <= na3274;

always @(posedge na3280)
   l358 <= na3280;

always @(posedge a3288)
   l360 <= a3288;

always @(posedge na3294)
   l362 <= na3294;

always @(posedge a3360)
   l364 <= a3360;

always @(posedge a3382)
   l366 <= a3382;

always @(posedge a3394)
   l368 <= a3394;

always @(posedge na3396)
   l370 <= na3396;

always @(posedge a3398)
   l372 <= a3398;

always @(posedge a3402)
   l374 <= a3402;

always @(posedge na3410)
   l376 <= na3410;

always @(posedge na3420)
   l378 <= na3420;

always @(posedge na1206)
   l380 <= na1206;

always @(posedge a3428)
   l382 <= a3428;

always @(posedge a1228)
   l384 <= a1228;

always @(posedge a1314)
   l386 <= a1314;

always @(posedge na3438)
   l388 <= na3438;

always @(posedge a1316)
   l390 <= a1316;

always @(posedge a3448)
   l392 <= a3448;

always @(posedge a3452)
   l394 <= a3452;

always @(posedge a3456)
   l396 <= a3456;

always @(posedge na3460)
   l398 <= na3460;

always @(posedge na3486)
   l400 <= na3486;

always @(posedge na3498)
   l402 <= na3498;

always @(posedge a1230)
   l404 <= a1230;

always @(posedge a3510)
   l406 <= a3510;

always @(posedge na3518)
   l408 <= na3518;

always @(posedge a3538)
   l410 <= a3538;

always @(posedge a3546)
   l412 <= a3546;

always @(posedge a3556)
   l414 <= a3556;

always @(posedge na2666)
   l416 <= na2666;

always @(posedge a3560)
   l418 <= a3560;

always @(posedge a3562)
   l420 <= a3562;

always @(posedge na3566)
   l422 <= na3566;

always @(posedge a3568)
   l424 <= a3568;

always @(posedge na3606)
   l426 <= na3606;

always @(posedge a3608)
   l428 <= a3608;

always @(posedge a3612)
   l430 <= a3612;

always @(posedge na3634)
   l432 <= na3634;

always @(posedge a3664)
   l434 <= a3664;

always @(posedge na3734)
   l436 <= na3734;

always @(posedge na3770)
   l438 <= na3770;

always @(posedge a3794)
   l440 <= a3794;

always @(posedge na3820)
   l442 <= na3820;

always @(posedge a3824)
   l444 <= a3824;

always @(posedge a3826)
   l446 <= a3826;

always @(posedge na3836)
   l448 <= na3836;

always @(posedge a3842)
   l450 <= a3842;

always @(posedge a3848)
   l452 <= a3848;

always @(posedge a3854)
   l454 <= a3854;

always @(posedge a3860)
   l456 <= a3860;

always @(posedge a3866)
   l458 <= a3866;

always @(posedge a3872)
   l460 <= a3872;

always @(posedge a3878)
   l462 <= a3878;

always @(posedge a3884)
   l464 <= a3884;

always @(posedge a3890)
   l466 <= a3890;

always @(posedge a3896)
   l468 <= a3896;

always @(posedge a3900)
   l470 <= a3900;

always @(posedge a1384)
   l472 <= a1384;

always @(posedge a1418)
   l474 <= a1418;

always @(posedge a3902)
   l476 <= a3902;

always @(posedge a3930)
   l478 <= a3930;

always @(posedge na1472)
   l480 <= na1472;

always @(posedge l830)
   l482 <= l830;

always @(posedge na3936)
   l484 <= na3936;

always @(posedge a3982)
   l486 <= a3982;

always @(posedge na1496)
   l488 <= na1496;

always @(posedge na4108)
   l490 <= na4108;

always @(posedge na4128)
   l492 <= na4128;

always @(posedge na4134)
   l494 <= na4134;

always @(posedge na4140)
   l496 <= na4140;

always @(posedge na4146)
   l498 <= na4146;

always @(posedge a4158)
   l500 <= a4158;

always @(posedge na4174)
   l502 <= na4174;

always @(posedge na4180)
   l504 <= na4180;

always @(posedge na4186)
   l506 <= na4186;

always @(posedge na4192)
   l508 <= na4192;

always @(posedge na4202)
   l510 <= na4202;

always @(posedge na4224)
   l512 <= na4224;

always @(posedge na4238)
   l514 <= na4238;

always @(posedge na4244)
   l516 <= na4244;

always @(posedge na4250)
   l518 <= na4250;

always @(posedge na4256)
   l520 <= na4256;

always @(posedge na4262)
   l522 <= na4262;

always @(posedge na4290)
   l524 <= na4290;

always @(posedge na4304)
   l526 <= na4304;

always @(posedge na4310)
   l528 <= na4310;

always @(posedge na4316)
   l530 <= na4316;

always @(posedge na4322)
   l532 <= na4322;

always @(posedge a4330)
   l534 <= a4330;

always @(posedge na4348)
   l536 <= na4348;

always @(posedge na4356)
   l538 <= na4356;

always @(posedge a4390)
   l540 <= a4390;

always @(posedge na4404)
   l542 <= na4404;

always @(posedge na4418)
   l544 <= na4418;

always @(posedge a4432)
   l546 <= a4432;

always @(posedge na4438)
   l548 <= na4438;

always @(posedge a4442)
   l550 <= a4442;

always @(posedge a4446)
   l552 <= a4446;

always @(posedge a4450)
   l554 <= a4450;

always @(posedge a4454)
   l556 <= a4454;

always @(posedge a4458)
   l558 <= a4458;

always @(posedge a4462)
   l560 <= a4462;

always @(posedge a4466)
   l562 <= a4466;

always @(posedge a4470)
   l564 <= a4470;

always @(posedge a4474)
   l566 <= a4474;

always @(posedge a4478)
   l568 <= a4478;

always @(posedge na4480)
   l570 <= na4480;

always @(posedge a4486)
   l572 <= a4486;

always @(posedge a4492)
   l574 <= a4492;

always @(posedge a4498)
   l576 <= a4498;

always @(posedge na4504)
   l578 <= na4504;

always @(posedge a4514)
   l580 <= a4514;

always @(posedge a4520)
   l582 <= a4520;

always @(posedge a4526)
   l584 <= a4526;

always @(posedge na4534)
   l586 <= na4534;

always @(posedge na4548)
   l588 <= na4548;

always @(posedge na4556)
   l590 <= na4556;

always @(posedge na4564)
   l592 <= na4564;

always @(posedge na4574)
   l594 <= na4574;

always @(posedge na4580)
   l596 <= na4580;

always @(posedge na4586)
   l598 <= na4586;

always @(posedge na4592)
   l600 <= na4592;

always @(posedge na4602)
   l602 <= na4602;

always @(posedge na4608)
   l604 <= na4608;

always @(posedge na4614)
   l606 <= na4614;

always @(posedge na4622)
   l608 <= na4622;

always @(posedge na4630)
   l610 <= na4630;

always @(posedge na4636)
   l612 <= na4636;

always @(posedge na4648)
   l614 <= na4648;

always @(posedge na4654)
   l616 <= na4654;

always @(posedge na4660)
   l618 <= na4660;

always @(posedge na4666)
   l620 <= na4666;

always @(posedge na4672)
   l622 <= na4672;

always @(posedge na4678)
   l624 <= na4678;

always @(posedge na4684)
   l626 <= na4684;

always @(posedge na4690)
   l628 <= na4690;

always @(posedge na4696)
   l630 <= na4696;

always @(posedge na4702)
   l632 <= na4702;

always @(posedge na4710)
   l634 <= na4710;

always @(posedge na4716)
   l636 <= na4716;

always @(posedge na4722)
   l638 <= na4722;

always @(posedge na4728)
   l640 <= na4728;

always @(posedge na4734)
   l642 <= na4734;

always @(posedge na4740)
   l644 <= na4740;

always @(posedge na4746)
   l646 <= na4746;

always @(posedge na4752)
   l648 <= na4752;

always @(posedge na4758)
   l650 <= na4758;

always @(posedge na4764)
   l652 <= na4764;

always @(posedge na4770)
   l654 <= na4770;

always @(posedge na4778)
   l656 <= na4778;

always @(posedge na4784)
   l658 <= na4784;

always @(posedge na4790)
   l660 <= na4790;

always @(posedge na4796)
   l662 <= na4796;

always @(posedge na4802)
   l664 <= na4802;

always @(posedge na4808)
   l666 <= na4808;

always @(posedge na4814)
   l668 <= na4814;

always @(posedge na4820)
   l670 <= na4820;

always @(posedge na4826)
   l672 <= na4826;

always @(posedge na4832)
   l674 <= na4832;

always @(posedge na4838)
   l676 <= na4838;

always @(posedge na4844)
   l678 <= na4844;

always @(posedge na4850)
   l680 <= na4850;

always @(posedge na4856)
   l682 <= na4856;

always @(posedge na4862)
   l684 <= na4862;

always @(posedge na4868)
   l686 <= na4868;

always @(posedge na4874)
   l688 <= na4874;

always @(posedge na4880)
   l690 <= na4880;

always @(posedge na4886)
   l692 <= na4886;

always @(posedge na4892)
   l694 <= na4892;

always @(posedge na4898)
   l696 <= na4898;

always @(posedge na4904)
   l698 <= na4904;

always @(posedge na4910)
   l700 <= na4910;

always @(posedge na4916)
   l702 <= na4916;

always @(posedge na4922)
   l704 <= na4922;

always @(posedge na4928)
   l706 <= na4928;

always @(posedge na4934)
   l708 <= na4934;

always @(posedge na4940)
   l710 <= na4940;

always @(posedge na4946)
   l712 <= na4946;

always @(posedge na4952)
   l714 <= na4952;

always @(posedge na4958)
   l716 <= na4958;

always @(posedge na4964)
   l718 <= na4964;

always @(posedge na4970)
   l720 <= na4970;

always @(posedge na4976)
   l722 <= na4976;

always @(posedge na4982)
   l724 <= na4982;

always @(posedge na4988)
   l726 <= na4988;

always @(posedge na4994)
   l728 <= na4994;

always @(posedge na5000)
   l730 <= na5000;

always @(posedge na5006)
   l732 <= na5006;

always @(posedge na5012)
   l734 <= na5012;

always @(posedge na5018)
   l736 <= na5018;

always @(posedge na5024)
   l738 <= na5024;

always @(posedge na5030)
   l740 <= na5030;

always @(posedge na5036)
   l742 <= na5036;

always @(posedge na5042)
   l744 <= na5042;

always @(posedge na5048)
   l746 <= na5048;

always @(posedge na5054)
   l748 <= na5054;

always @(posedge na5060)
   l750 <= na5060;

always @(posedge na5066)
   l752 <= na5066;

always @(posedge na5072)
   l754 <= na5072;

always @(posedge na5078)
   l756 <= na5078;

always @(posedge na5084)
   l758 <= na5084;

always @(posedge na5090)
   l760 <= na5090;

always @(posedge na5096)
   l762 <= na5096;

always @(posedge na5102)
   l764 <= na5102;

always @(posedge na5108)
   l766 <= na5108;

always @(posedge na5114)
   l768 <= na5114;

always @(posedge na5120)
   l770 <= na5120;

always @(posedge na5126)
   l772 <= na5126;

always @(posedge na5132)
   l774 <= na5132;

always @(posedge na5138)
   l776 <= na5138;

always @(posedge na5144)
   l778 <= na5144;

always @(posedge na5150)
   l780 <= na5150;

always @(posedge na5156)
   l782 <= na5156;

always @(posedge na5162)
   l784 <= na5162;

always @(posedge na5168)
   l786 <= na5168;

always @(posedge na5174)
   l788 <= na5174;

always @(posedge na5180)
   l790 <= na5180;

always @(posedge na5186)
   l792 <= na5186;

always @(posedge na5192)
   l794 <= na5192;

always @(posedge na5198)
   l796 <= na5198;

always @(posedge na5204)
   l798 <= na5204;

always @(posedge na5210)
   l800 <= na5210;

always @(posedge na5216)
   l802 <= na5216;

always @(posedge na5222)
   l804 <= na5222;

always @(posedge na5228)
   l806 <= na5228;

always @(posedge na5234)
   l808 <= na5234;

always @(posedge na5240)
   l810 <= na5240;

always @(posedge na5244)
   l812 <= na5244;

always @(posedge a5250)
   l814 <= a5250;

always @(posedge na5262)
   l816 <= na5262;

always @(posedge na5274)
   l818 <= na5274;

always @(posedge na5286)
   l820 <= na5286;

always @(posedge a5296)
   l822 <= a5296;

always @(posedge a5298)
   l824 <= a5298;

always @(posedge a5300)
   l826 <= a5300;

always @(posedge na5308)
   l828 <= na5308;

always @(posedge a5310)
   l830 <= a5310;

always @(posedge a5312)
   l832 <= a5312;

always @(posedge na5316)
   l834 <= na5316;

always @(posedge na5320)
   l836 <= na5320;

always @(posedge a5322)
   l838 <= a5322;

always @(posedge a5326)
   l840 <= a5326;

always @(posedge na5330)
   l842 <= na5330;

always @(posedge a5332)
   l844 <= a5332;

always @(posedge a5340)
   l846 <= a5340;

always @(posedge a5346)
   l848 <= a5346;

always @(posedge a5352)
   l850 <= a5352;

always @(posedge a5362)
   l852 <= a5362;

always @(posedge na5414)
   l854 <= na5414;

always @(posedge a5424)
   l856 <= a5424;

always @(posedge na5442)
   l858 <= na5442;

always @(posedge a5444)
   l860 <= a5444;

always @(posedge a5450)
   l862 <= a5450;

always @(posedge na5456)
   l864 <= na5456;

always @(posedge a5464)
   l866 <= a5464;

always @(posedge a5472)
   l868 <= a5472;

always @(posedge a5480)
   l870 <= a5480;

always @(posedge a5492)
   l872 <= a5492;

always @(posedge a5500)
   l874 <= a5500;

always @(posedge a5510)
   l876 <= a5510;

always @(posedge a5518)
   l878 <= a5518;

always @(posedge a5526)
   l880 <= a5526;

always @(posedge a5534)
   l882 <= a5534;

always @(posedge a5540)
   l884 <= a5540;

always @(posedge a5546)
   l886 <= a5546;

always @(posedge a5552)
   l888 <= a5552;

always @(posedge a5558)
   l890 <= a5558;

always @(posedge a5564)
   l892 <= a5564;

always @(posedge a5570)
   l894 <= a5570;

always @(posedge a5578)
   l896 <= a5578;

always @(posedge a5584)
   l898 <= a5584;

always @(posedge a5590)
   l900 <= a5590;

always @(posedge a5596)
   l902 <= a5596;

always @(posedge a5602)
   l904 <= a5602;

always @(posedge a5608)
   l906 <= a5608;

always @(posedge a5614)
   l908 <= a5614;

always @(posedge a5622)
   l910 <= a5622;

always @(posedge a5628)
   l912 <= a5628;

always @(posedge a5634)
   l914 <= a5634;

always @(posedge a5640)
   l916 <= a5640;

always @(posedge a5646)
   l918 <= a5646;

always @(posedge a5652)
   l920 <= a5652;

always @(posedge a5660)
   l922 <= a5660;

always @(posedge a5666)
   l924 <= a5666;

always @(posedge a5672)
   l926 <= a5672;

always @(posedge a5678)
   l928 <= a5678;

always @(posedge a5684)
   l930 <= a5684;

always @(posedge a5690)
   l932 <= a5690;

always @(posedge a5696)
   l934 <= a5696;

always @(posedge a5704)
   l936 <= a5704;

always @(posedge a5710)
   l938 <= a5710;

always @(posedge a5716)
   l940 <= a5716;

always @(posedge a5722)
   l942 <= a5722;

always @(posedge a5728)
   l944 <= a5728;

always @(posedge a5734)
   l946 <= a5734;

always @(posedge a5740)
   l948 <= a5740;

always @(posedge a5748)
   l950 <= a5748;

always @(posedge a5754)
   l952 <= a5754;

always @(posedge a5760)
   l954 <= a5760;

always @(posedge a5766)
   l956 <= a5766;

always @(posedge a5772)
   l958 <= a5772;

always @(posedge a5778)
   l960 <= a5778;

always @(posedge a5784)
   l962 <= a5784;

always @(posedge a5792)
   l964 <= a5792;

always @(posedge a5798)
   l966 <= a5798;

always @(posedge a5804)
   l968 <= a5804;

always @(posedge a5810)
   l970 <= a5810;

always @(posedge a5816)
   l972 <= a5816;

always @(posedge a5822)
   l974 <= a5822;

always @(posedge a5828)
   l976 <= a5828;

always @(posedge na5830)
   l978 <= na5830;

always @(posedge a5834)
   l980 <= a5834;

always @(posedge a5888)
   l982 <= a5888;

always @(posedge a5918)
   l984 <= a5918;

always @(posedge a5948)
   l986 <= a5948;

always @(posedge a5978)
   l988 <= a5978;

always @(posedge a6008)
   l990 <= a6008;

always @(posedge na6102)
   l992 <= na6102;

always @(posedge a6106)
   l994 <= a6106;

always @(posedge a6110)
   l996 <= a6110;

always @(posedge a6112)
   l998 <= a6112;

always @(posedge a6114)
   l1000 <= a6114;

always @(posedge a6116)
   l1002 <= a6116;

always @(posedge na6138)
   l1004 <= na6138;

always @(posedge na6148)
   l1006 <= na6148;


assign na2642 = ~a2642;
assign a2694 = ~a2692 & ~a2598;
assign na2694 = ~a2694;
assign na2622 = ~a2622;
assign a2582 = ~a2580 & ~a2578;
assign na2576 = ~a2576;
assign na2570 = ~a2570;
assign na2564 = ~a2564;
assign na2558 = ~a2558;
assign na2616 = ~a2616;
assign na2610 = ~a2610;
assign na2698 = ~a2698;
assign na2632 = ~a2632;
assign na2604 = ~a2604;
assign c1 = 1;
assign a2546 = l274 & i42;
assign a2704 = ~a2702 & ~a2700;
assign a2710 = ~a2708 & ~a2706;
assign a2712 = l996 & ~l292;
assign a2774 = ~a2772 & ~a2770;
assign a2778 = ~a2776 & ~a1012;
assign na2780 = ~a2780;
assign na2816 = ~a2816;
assign a2838 = ~a2836 & ~a2832;
assign a2842 = ~a2840 & ~a1026;
assign na2846 = ~a2846;
assign na2850 = ~a2850;
assign na2856 = ~a2856;
assign na2862 = ~a2862;
assign na2868 = ~a2868;
assign na2874 = ~a2874;
assign na2880 = ~a2880;
assign na2886 = ~a2886;
assign na2892 = ~a2892;
assign na2898 = ~a2898;
assign na2904 = ~a2904;
assign na2908 = ~a2908;
assign a2910 = ~a2906 & a2780;
assign a2916 = ~a2914 & l854;
assign a3060 = ~a3058 & ~a3046;
assign a3080 = ~a3078 & ~a3062;
assign a3200 = ~a3198 & ~a3156;
assign na3230 = ~a3230;
assign a3232 = a2550 & ~a2546;
assign na3238 = ~a3238;
assign na3244 = ~a3244;
assign na3250 = ~a3250;
assign na3256 = ~a3256;
assign na3262 = ~a3262;
assign na3268 = ~a3268;
assign na3274 = ~a3274;
assign na3280 = ~a3280;
assign a3288 = ~a3286 & ~a3284;
assign na3294 = ~a3294;
assign a3360 = ~a3358 & ~a3336;
assign a3382 = ~a3380 & ~a3378;
assign a3394 = ~a3392 & ~a3384;
assign na3396 = ~a3396;
assign a3398 = a3396 & a3360;
assign a3402 = ~a3400 & a3396;
assign na3410 = ~a3410;
assign na3420 = ~a3420;
assign na1206 = ~a1206;
assign a3428 = ~a3426 & ~a1262;
assign a1228 = ~a1226 & ~a1208;
assign a1314 = ~a1312 & ~a1310;
assign na3438 = ~a3438;
assign a1316 = a1314 & a1298;
assign a3448 = ~a3446 & ~a3442;
assign a3452 = ~a3450 & ~a3416;
assign a3456 = a3454 & ~a3394;
assign na3460 = ~a3460;
assign na3486 = ~a3486;
assign na3498 = ~a3498;
assign a1230 = a1228 & ~a1206;
assign a3510 = ~a3508 & a3500;
assign na3518 = ~a3518;
assign a3538 = ~a3536 & l370;
assign a3546 = ~a3544 & l370;
assign a3556 = ~a3554 & ~a2652;
assign na2666 = ~a2666;
assign a3560 = ~a3558 & ~a3282;
assign a3562 = a3404 & l422;
assign na3566 = ~a3566;
assign a3568 = a3462 & ~a1314;
assign na3606 = ~a3606;
assign a3608 = l430 & l302;
assign a3612 = ~a3610 & ~a3608;
assign na3634 = ~a3634;
assign a3664 = ~a3662 & ~a3636;
assign na3734 = ~a3734;
assign na3770 = ~a3770;
assign a3794 = ~a3792 & ~a3772;
assign na3820 = ~a3820;
assign a3824 = a3822 & ~a1250;
assign a3826 = ~a2652 & ~a1254;
assign na3836 = ~a3836;
assign a3842 = a3840 & ~a1010;
assign a3848 = a3846 & ~a1278;
assign a3854 = a3852 & ~a1280;
assign a3860 = a3858 & ~a1282;
assign a3866 = a3864 & ~a1284;
assign a3872 = a3870 & ~a1286;
assign a3878 = a3876 & ~a1288;
assign a3884 = a3882 & ~a1290;
assign a3890 = a3888 & ~a1292;
assign a3896 = a3894 & ~a1294;
assign a3900 = ~a3898 & ~a1010;
assign a1384 = ~a1382 & a1338;
assign a1418 = a1416 & ~a1412;
assign a3902 = ~l426 & l406;
assign a3930 = ~a3928 & ~a1444;
assign na1472 = ~a1472;
assign na3936 = ~a3936;
assign a3982 = ~a3980 & ~a2552;
assign na1496 = ~a1496;
assign na4108 = ~a4108;
assign na4128 = ~a4128;
assign na4134 = ~a4134;
assign na4140 = ~a4140;
assign na4146 = ~a4146;
assign a4158 = ~a4156 & ~a4148;
assign na4174 = ~a4174;
assign na4180 = ~a4180;
assign na4186 = ~a4186;
assign na4192 = ~a4192;
assign na4202 = ~a4202;
assign na4224 = ~a4224;
assign na4238 = ~a4238;
assign na4244 = ~a4244;
assign na4250 = ~a4250;
assign na4256 = ~a4256;
assign na4262 = ~a4262;
assign na4290 = ~a4290;
assign na4304 = ~a4304;
assign na4310 = ~a4310;
assign na4316 = ~a4316;
assign na4322 = ~a4322;
assign a4330 = ~a4328 & ~a4274;
assign na4348 = ~a4348;
assign na4356 = ~a4356;
assign a4390 = ~a4388 & ~a4374;
assign na4404 = ~a4404;
assign na4418 = ~a4418;
assign a4432 = ~a4430 & ~a4428;
assign na4438 = ~a4438;
assign a4442 = ~a4440 & ~a1682;
assign a4446 = ~a4444 & ~a1684;
assign a4450 = ~a4448 & ~a1686;
assign a4454 = ~a4452 & ~a1688;
assign a4458 = ~a4456 & ~a1690;
assign a4462 = ~a4460 & ~a1692;
assign a4466 = ~a4464 & ~a1694;
assign a4470 = ~a4468 & ~a1696;
assign a4474 = ~a4472 & ~a1698;
assign a4478 = ~a4476 & ~a1700;
assign na4480 = ~a4480;
assign a4486 = ~a4484 & ~a4482;
assign a4492 = ~a4490 & ~a4488;
assign a4498 = ~a4496 & ~a4494;
assign na4504 = ~a4504;
assign a4514 = ~a4512 & ~a4510;
assign a4520 = ~a4518 & ~a4516;
assign a4526 = ~a4524 & ~a4522;
assign na4534 = ~a4534;
assign na4548 = ~a4548;
assign na4556 = ~a4556;
assign na4564 = ~a4564;
assign na4574 = ~a4574;
assign na4580 = ~a4580;
assign na4586 = ~a4586;
assign na4592 = ~a4592;
assign na4602 = ~a4602;
assign na4608 = ~a4608;
assign na4614 = ~a4614;
assign na4622 = ~a4622;
assign na4630 = ~a4630;
assign na4636 = ~a4636;
assign na4648 = ~a4648;
assign na4654 = ~a4654;
assign na4660 = ~a4660;
assign na4666 = ~a4666;
assign na4672 = ~a4672;
assign na4678 = ~a4678;
assign na4684 = ~a4684;
assign na4690 = ~a4690;
assign na4696 = ~a4696;
assign na4702 = ~a4702;
assign na4710 = ~a4710;
assign na4716 = ~a4716;
assign na4722 = ~a4722;
assign na4728 = ~a4728;
assign na4734 = ~a4734;
assign na4740 = ~a4740;
assign na4746 = ~a4746;
assign na4752 = ~a4752;
assign na4758 = ~a4758;
assign na4764 = ~a4764;
assign na4770 = ~a4770;
assign na4778 = ~a4778;
assign na4784 = ~a4784;
assign na4790 = ~a4790;
assign na4796 = ~a4796;
assign na4802 = ~a4802;
assign na4808 = ~a4808;
assign na4814 = ~a4814;
assign na4820 = ~a4820;
assign na4826 = ~a4826;
assign na4832 = ~a4832;
assign na4838 = ~a4838;
assign na4844 = ~a4844;
assign na4850 = ~a4850;
assign na4856 = ~a4856;
assign na4862 = ~a4862;
assign na4868 = ~a4868;
assign na4874 = ~a4874;
assign na4880 = ~a4880;
assign na4886 = ~a4886;
assign na4892 = ~a4892;
assign na4898 = ~a4898;
assign na4904 = ~a4904;
assign na4910 = ~a4910;
assign na4916 = ~a4916;
assign na4922 = ~a4922;
assign na4928 = ~a4928;
assign na4934 = ~a4934;
assign na4940 = ~a4940;
assign na4946 = ~a4946;
assign na4952 = ~a4952;
assign na4958 = ~a4958;
assign na4964 = ~a4964;
assign na4970 = ~a4970;
assign na4976 = ~a4976;
assign na4982 = ~a4982;
assign na4988 = ~a4988;
assign na4994 = ~a4994;
assign na5000 = ~a5000;
assign na5006 = ~a5006;
assign na5012 = ~a5012;
assign na5018 = ~a5018;
assign na5024 = ~a5024;
assign na5030 = ~a5030;
assign na5036 = ~a5036;
assign na5042 = ~a5042;
assign na5048 = ~a5048;
assign na5054 = ~a5054;
assign na5060 = ~a5060;
assign na5066 = ~a5066;
assign na5072 = ~a5072;
assign na5078 = ~a5078;
assign na5084 = ~a5084;
assign na5090 = ~a5090;
assign na5096 = ~a5096;
assign na5102 = ~a5102;
assign na5108 = ~a5108;
assign na5114 = ~a5114;
assign na5120 = ~a5120;
assign na5126 = ~a5126;
assign na5132 = ~a5132;
assign na5138 = ~a5138;
assign na5144 = ~a5144;
assign na5150 = ~a5150;
assign na5156 = ~a5156;
assign na5162 = ~a5162;
assign na5168 = ~a5168;
assign na5174 = ~a5174;
assign na5180 = ~a5180;
assign na5186 = ~a5186;
assign na5192 = ~a5192;
assign na5198 = ~a5198;
assign na5204 = ~a5204;
assign na5210 = ~a5210;
assign na5216 = ~a5216;
assign na5222 = ~a5222;
assign na5228 = ~a5228;
assign na5234 = ~a5234;
assign na5240 = ~a5240;
assign na5244 = ~a5244;
assign a5250 = ~a5248 & ~a5246;
assign na5262 = ~a5262;
assign na5274 = ~a5274;
assign na5286 = ~a5286;
assign a5296 = ~a5294 & ~a5290;
assign a5298 = a3824 & a2664;
assign a5300 = l980 & ~l826;
assign na5308 = ~a5308;
assign a5310 = ~a3606 & ~l426;
assign a5312 = ~a2638 & ~a2584;
assign na5316 = ~a5316;
assign na5320 = ~a5320;
assign a5322 = ~a2588 & a2558;
assign a5326 = ~a5324 & ~a2624;
assign na5330 = ~a5330;
assign a5332 = ~a2634 & a2604;
assign a5340 = a5338 & ~a5334;
assign a5346 = ~a5344 & ~a5342;
assign a5352 = ~a5350 & ~a5348;
assign a5362 = ~a5360 & ~a5358;
assign na5414 = ~a5414;
assign a5424 = a5422 & ~a5418;
assign na5442 = ~a5442;
assign a5444 = ~a5436 & ~a2912;
assign a5450 = ~a5448 & ~a5446;
assign na5456 = ~a5456;
assign a5464 = ~a5462 & ~a5460;
assign a5472 = ~a5470 & ~a5468;
assign a5480 = ~a5478 & ~a5476;
assign a5492 = ~a5490 & ~a5488;
assign a5500 = ~a5498 & ~a5496;
assign a5510 = ~a5508 & ~a5506;
assign a5518 = ~a5516 & ~a5514;
assign a5526 = ~a5524 & ~a5522;
assign a5534 = ~a5532 & ~a5530;
assign a5540 = ~a5538 & ~a5536;
assign a5546 = ~a5544 & ~a5542;
assign a5552 = ~a5550 & ~a5548;
assign a5558 = ~a5556 & ~a5554;
assign a5564 = ~a5562 & ~a5560;
assign a5570 = ~a5568 & ~a5566;
assign a5578 = ~a5576 & ~a5574;
assign a5584 = ~a5582 & ~a5580;
assign a5590 = ~a5588 & ~a5586;
assign a5596 = ~a5594 & ~a5592;
assign a5602 = ~a5600 & ~a5598;
assign a5608 = ~a5606 & ~a5604;
assign a5614 = ~a5612 & ~a5610;
assign a5622 = ~a5620 & ~a5618;
assign a5628 = ~a5626 & ~a5624;
assign a5634 = ~a5632 & ~a5630;
assign a5640 = ~a5638 & ~a5636;
assign a5646 = ~a5644 & ~a5642;
assign a5652 = ~a5650 & ~a5648;
assign a5660 = ~a5658 & ~a5656;
assign a5666 = ~a5664 & ~a5662;
assign a5672 = ~a5670 & ~a5668;
assign a5678 = ~a5676 & ~a5674;
assign a5684 = ~a5682 & ~a5680;
assign a5690 = ~a5688 & ~a5686;
assign a5696 = ~a5694 & ~a5692;
assign a5704 = ~a5702 & ~a5700;
assign a5710 = ~a5708 & ~a5706;
assign a5716 = ~a5714 & ~a5712;
assign a5722 = ~a5720 & ~a5718;
assign a5728 = ~a5726 & ~a5724;
assign a5734 = ~a5732 & ~a5730;
assign a5740 = ~a5738 & ~a5736;
assign a5748 = ~a5746 & ~a5744;
assign a5754 = ~a5752 & ~a5750;
assign a5760 = ~a5758 & ~a5756;
assign a5766 = ~a5764 & ~a5762;
assign a5772 = ~a5770 & ~a5768;
assign a5778 = ~a5776 & ~a5774;
assign a5784 = ~a5782 & ~a5780;
assign a5792 = ~a5790 & ~a5788;
assign a5798 = ~a5796 & ~a5794;
assign a5804 = ~a5802 & ~a5800;
assign a5810 = ~a5808 & ~a5806;
assign a5816 = ~a5814 & ~a5812;
assign a5822 = ~a5820 & ~a5818;
assign a5828 = ~a5826 & ~a5824;
assign na5830 = ~a5830;
assign a5834 = a5832 & ~a5416;
assign a5888 = a5886 & a5862;
assign a5918 = a5916 & a5902;
assign a5948 = a5946 & a5932;
assign a5978 = a5976 & a5962;
assign a6008 = a6006 & a5992;
assign na6102 = ~a6102;
assign a6106 = a6104 & ~l1006;
assign a6110 = a6108 & a2816;
assign a6112 = a6110 & ~l1002;
assign a6114 = a6112 & l998;
assign a6116 = a6114 & ~a2712;
assign na6138 = ~a6138;
assign na6148 = ~a6148;
assign a1008 = l368 & l366;
assign a1010 = a1008 & l364;
assign a1012 = ~a1010 & ~l296;
assign a1014 = l300 & l294;
assign a1016 = a1014 & l298;
assign a1018 = ~a1016 & ~l328;
assign a1020 = ~a1018 & l340;
assign a1022 = ~a1020 & ~l996;
assign a1024 = ~a1022 & a1012;
assign a1026 = l432 & l304;
assign a1028 = a1026 & l306;
assign a1030 = a1028 & l308;
assign a1032 = a1030 & l374;
assign a1034 = l432 & ~l304;
assign a1036 = a1034 & l306;
assign a1038 = a1036 & l308;
assign a1040 = a1038 & l374;
assign a1042 = a1026 & ~l306;
assign a1044 = a1042 & l308;
assign a1046 = a1044 & l374;
assign a1048 = a1034 & ~l306;
assign a1050 = a1048 & l308;
assign a1052 = a1050 & l374;
assign a1054 = a1028 & ~l308;
assign a1056 = a1054 & l374;
assign a1058 = a1036 & ~l308;
assign a1060 = a1058 & l374;
assign a1062 = a1042 & ~l308;
assign a1064 = a1062 & l374;
assign a1066 = a1048 & ~l308;
assign a1068 = a1066 & l374;
assign a1070 = l372 & l282;
assign a1072 = l426 & l408;
assign a1074 = a1072 & ~l422;
assign a1076 = a1074 & ~a1070;
assign a1078 = l828 & ~l376;
assign a1080 = ~a1078 & l378;
assign a1082 = l378 & l372;
assign a1084 = l386 & ~l384;
assign a1086 = a1084 & l380;
assign a1088 = ~l402 & ~l400;
assign a1090 = ~l382 & l276;
assign a1092 = a1090 & l278;
assign a1094 = a1092 & a1088;
assign a1096 = a1094 & a1086;
assign a1098 = ~l402 & l400;
assign a1100 = a1098 & l382;
assign a1102 = l408 & l388;
assign a1104 = a1102 & a1094;
assign a1106 = a1102 & ~a1092;
assign a1108 = l274 & i54;
assign a1110 = l274 & i60;
assign a1112 = l274 & i58;
assign a1114 = a1112 & ~a1110;
assign a1116 = a1114 & ~i56;
assign a1118 = a1116 & a1108;
assign a1120 = ~l402 & l388;
assign a1122 = ~a1120 & l408;
assign a1124 = a1122 & a1118;
assign a1126 = ~a1124 & ~a1094;
assign a1128 = ~a1126 & l404;
assign a1130 = ~l386 & ~l384;
assign a1132 = a1130 & l380;
assign a1134 = a1090 & a1086;
assign a1136 = ~a1134 & ~a1132;
assign a1138 = a1136 & ~a1128;
assign a1140 = a1138 & l380;
assign a1142 = a1090 & ~l278;
assign a1144 = a1142 & a1088;
assign a1146 = l274 & i56;
assign a1148 = ~a1146 & a1108;
assign a1150 = ~l278 & l276;
assign a1152 = a1150 & ~a1098;
assign a1154 = a1152 & a1148;
assign a1156 = ~a1154 & ~a1144;
assign a1158 = ~a1156 & l390;
assign a1160 = a1130 & ~l380;
assign a1162 = a1160 & l396;
assign a1164 = ~a1162 & ~a1158;
assign a1166 = a1164 & a1138;
assign a1168 = l274 & ~i50;
assign a1170 = a1168 & i48;
assign a1172 = ~a1170 & ~l386;
assign a1174 = l384 & ~l380;
assign a1176 = a1174 & ~a1172;
assign a1178 = ~a1176 & a1166;
assign a1180 = a1142 & l402;
assign a1182 = a1180 & a1148;
assign a1184 = a1182 & l390;
assign a1186 = a1172 & ~l384;
assign a1188 = ~a1142 & a1086;
assign a1190 = a1102 & l404;
assign a1192 = l424 & l278;
assign a1194 = ~a1192 & ~a1160;
assign a1196 = a1194 & ~a1190;
assign a1198 = a1196 & ~a1188;
assign a1200 = a1198 & ~a1186;
assign a1202 = a1200 & ~a1184;
assign a1204 = ~a1202 & ~a1178;
assign a1206 = ~a1204 & ~a1140;
assign a1208 = a1166 & ~l384;
assign a1210 = ~a1182 & l390;
assign a1212 = a1170 & a1132;
assign a1214 = ~a1150 & l424;
assign a1216 = ~a1102 & l404;
assign a1218 = ~a1216 & ~a1214;
assign a1220 = a1218 & ~a1212;
assign a1222 = a1220 & ~a1188;
assign a1224 = a1222 & ~a1210;
assign a1226 = a1224 & ~a1178;
assign a1232 = a1230 & l278;
assign a1234 = a1232 & a1098;
assign a1236 = a1234 & ~a1102;
assign a1238 = ~l414 & ~l412;
assign a1240 = a1238 & ~l410;
assign a1242 = a1078 & l416;
assign a1244 = a1242 & ~a1240;
assign a1246 = a1142 & ~l444;
assign a1248 = a1246 & ~a1244;
assign a1250 = a1244 & l444;
assign a1252 = a1250 & l446;
assign a1254 = ~a1250 & ~l446;
assign a1256 = a1254 & l824;
assign a1258 = ~a1256 & ~a1252;
assign a1260 = ~l368 & l366;
assign a1262 = a1260 & l378;
assign a1264 = a1262 & ~l364;
assign a1266 = a1264 & a1240;
assign a1268 = l824 & l446;
assign a1270 = ~a1268 & a1266;
assign a1272 = a1268 & ~a1266;
assign a1274 = ~a1272 & ~a1270;
assign a1276 = l450 & l448;
assign a1278 = a1276 & l452;
assign a1280 = a1278 & l454;
assign a1282 = a1280 & l456;
assign a1284 = a1282 & l458;
assign a1286 = a1284 & l460;
assign a1288 = a1286 & l462;
assign a1290 = a1288 & l464;
assign a1292 = a1290 & l466;
assign a1294 = a1292 & l468;
assign a1296 = a1294 & l470;
assign a1298 = ~a1228 & a1206;
assign a1300 = a1142 & a1086;
assign a1302 = a1150 & l424;
assign a1304 = ~l404 & ~l390;
assign a1306 = a1304 & ~a1302;
assign a1308 = a1306 & ~a1300;
assign a1310 = a1308 & ~a1178;
assign a1312 = a1178 & ~l386;
assign a1318 = ~a1148 & a1144;
assign a1320 = a1318 & a1316;
assign a1322 = l830 & l406;
assign a1324 = ~a1146 & ~a1108;
assign a1326 = ~a1112 & ~a1110;
assign a1328 = a1326 & a1324;
assign a1330 = ~i8 & ~i6;
assign a1332 = a1330 & ~a1114;
assign a1334 = ~a1332 & ~a1328;
assign a1336 = ~l426 & ~l406;
assign a1338 = ~a1336 & ~l830;
assign a1340 = ~l478 & l472;
assign a1342 = ~l480 & ~l474;
assign a1344 = a1342 & a1340;
assign a1346 = l480 & l474;
assign a1348 = a1346 & ~l472;
assign a1350 = ~a1348 & ~a1344;
assign a1352 = ~a1350 & ~a1338;
assign a1354 = a1108 & l406;
assign a1356 = ~a1354 & a1116;
assign a1358 = ~a1356 & a1352;
assign a1360 = a1358 & a1334;
assign a1362 = l474 & ~l472;
assign a1364 = a1362 & ~l480;
assign a1366 = ~a1364 & ~l482;
assign a1368 = ~a1366 & ~a1338;
assign a1370 = ~a1346 & a1340;
assign a1372 = a1370 & ~a1342;
assign a1374 = a1372 & a1356;
assign a1376 = ~a1338 & ~l476;
assign a1378 = a1376 & a1374;
assign a1380 = ~a1330 & a1328;
assign a1382 = a1380 & ~a1366;
assign a1386 = a1342 & ~l472;
assign a1388 = a1386 & a1384;
assign a1390 = ~a1356 & a1338;
assign a1392 = a1390 & l476;
assign a1394 = l478 & ~l474;
assign a1396 = a1394 & ~a1392;
assign a1398 = a1350 & a1338;
assign a1400 = a1398 & ~a1374;
assign a1402 = a1400 & ~a1396;
assign a1404 = ~a1402 & ~a1366;
assign a1406 = ~a1390 & a1334;
assign a1408 = ~a1380 & ~a1350;
assign a1410 = a1408 & ~a1406;
assign a1412 = ~a1410 & ~a1402;
assign a1414 = a1406 & ~a1366;
assign a1416 = ~a1414 & ~a1386;
assign a1420 = a1382 & a1338;
assign a1422 = a1420 & ~a1418;
assign a1424 = a1418 & ~a1338;
assign a1426 = ~a1424 & ~a1422;
assign a1428 = ~a1392 & ~l830;
assign a1430 = a1428 & ~a1116;
assign a1432 = a1354 & a1116;
assign a1434 = ~a1432 & ~a1430;
assign a1436 = ~a1434 & ~l476;
assign a1438 = a1336 & l476;
assign a1440 = ~a1438 & a1372;
assign a1442 = a1440 & ~a1436;
assign a1444 = a1346 & a1340;
assign a1446 = a1444 & ~a1336;
assign a1448 = ~a1446 & a1428;
assign a1450 = a1448 & ~a1442;
assign a1452 = ~a1362 & ~a1344;
assign a1454 = a1452 & ~a1450;
assign a1456 = ~a1434 & a1334;
assign a1458 = ~a1456 & a1364;
assign a1460 = a1434 & ~a1328;
assign a1462 = ~a1460 & ~a1332;
assign a1464 = l480 & ~l472;
assign a1466 = ~a1464 & ~a1344;
assign a1468 = ~a1466 & ~a1462;
assign a1470 = ~a1468 & ~a1458;
assign a1472 = a1470 & ~a1454;
assign a1474 = a1386 & ~l830;
assign a1476 = a1474 & ~a1472;
assign a1478 = a1472 & l830;
assign a1480 = ~a1472 & a1336;
assign a1482 = ~a1480 & ~a1478;
assign a1484 = a1336 & l484;
assign a1486 = a1484 & a1326;
assign a1488 = a1336 & ~l476;
assign a1490 = ~a1488 & a1474;
assign a1492 = a1488 & ~a1474;
assign a1494 = ~a1492 & ~a1490;
assign a1496 = ~l438 & ~l436;
assign a1498 = ~l442 & ~l440;
assign a1500 = a1498 & ~l340;
assign a1502 = ~a1500 & ~a1496;
assign a1504 = a1500 & a1496;
assign a1506 = ~a1504 & ~a1502;
assign a1508 = ~l526 & i30;
assign a1510 = l528 & ~i34;
assign a1512 = ~a1510 & ~a1508;
assign a1514 = l526 & ~i30;
assign a1516 = ~l528 & i34;
assign a1518 = ~a1516 & ~a1514;
assign a1520 = a1518 & a1512;
assign a1522 = l274 & i38;
assign a1524 = ~a1522 & l530;
assign a1526 = a1522 & ~l530;
assign a1528 = ~a1526 & ~a1524;
assign a1530 = a1528 & a1520;
assign a1532 = ~i46 & ~i32;
assign a1534 = ~i40 & ~i36;
assign a1536 = a1534 & a1532;
assign a1538 = ~a1536 & l274;
assign a1540 = l274 & i44;
assign a1542 = a1540 & l532;
assign a1544 = ~a1540 & ~l532;
assign a1546 = ~a1544 & ~a1542;
assign a1548 = ~a1546 & ~a1538;
assign a1550 = a1548 & a1530;
assign a1552 = a1550 & l534;
assign a1554 = ~l492 & i30;
assign a1556 = l494 & ~i34;
assign a1558 = ~a1556 & ~a1554;
assign a1560 = l492 & ~i30;
assign a1562 = ~l494 & i34;
assign a1564 = ~a1562 & ~a1560;
assign a1566 = a1564 & a1558;
assign a1568 = ~a1540 & l498;
assign a1570 = a1540 & ~l498;
assign a1572 = ~a1570 & ~a1568;
assign a1574 = a1572 & a1566;
assign a1576 = a1522 & l496;
assign a1578 = ~a1522 & ~l496;
assign a1580 = ~a1578 & ~a1576;
assign a1582 = ~a1580 & ~a1538;
assign a1584 = a1582 & a1574;
assign a1586 = a1584 & l500;
assign a1588 = a1586 & a1552;
assign a1590 = ~l502 & i30;
assign a1592 = l504 & ~i34;
assign a1594 = ~a1592 & ~a1590;
assign a1596 = l502 & ~i30;
assign a1598 = ~l504 & i34;
assign a1600 = ~a1598 & ~a1596;
assign a1602 = a1600 & a1594;
assign a1604 = ~a1540 & l508;
assign a1606 = a1540 & ~l508;
assign a1608 = ~a1606 & ~a1604;
assign a1610 = a1608 & a1602;
assign a1612 = a1522 & l506;
assign a1614 = ~a1522 & ~l506;
assign a1616 = ~a1614 & ~a1612;
assign a1618 = ~a1616 & ~a1538;
assign a1620 = a1618 & a1610;
assign a1622 = a1620 & l510;
assign a1624 = ~a1622 & ~a1586;
assign a1626 = ~l514 & i30;
assign a1628 = l516 & ~i34;
assign a1630 = ~a1628 & ~a1626;
assign a1632 = l514 & ~i30;
assign a1634 = ~l516 & i34;
assign a1636 = ~a1634 & ~a1632;
assign a1638 = a1636 & a1630;
assign a1640 = ~a1540 & l520;
assign a1642 = a1540 & ~l520;
assign a1644 = ~a1642 & ~a1640;
assign a1646 = a1644 & a1638;
assign a1648 = a1522 & l518;
assign a1650 = ~a1522 & ~l518;
assign a1652 = ~a1650 & ~a1648;
assign a1654 = ~a1652 & ~a1538;
assign a1656 = a1654 & a1646;
assign a1658 = a1656 & l522;
assign a1660 = a1658 & ~a1624;
assign a1662 = ~a1658 & a1624;
assign a1664 = ~a1662 & a1552;
assign a1666 = ~a1622 & ~a1552;
assign a1668 = ~a1666 & a1658;
assign a1670 = ~a1496 & ~l488;
assign a1672 = ~l548 & ~l540;
assign a1674 = a1672 & ~l542;
assign a1676 = ~l546 & ~l544;
assign a1678 = a1676 & a1674;
assign a1680 = a1678 & ~a1670;
assign a1682 = ~a1680 & l550;
assign a1684 = a1682 & l552;
assign a1686 = a1684 & l554;
assign a1688 = a1686 & l556;
assign a1690 = a1688 & l558;
assign a1692 = a1690 & l560;
assign a1694 = a1692 & l562;
assign a1696 = a1694 & l564;
assign a1698 = a1696 & l566;
assign a1700 = a1698 & l568;
assign a1702 = a1700 & l570;
assign a1704 = ~l574 & ~l572;
assign a1706 = l578 & ~l576;
assign a1708 = a1706 & a1704;
assign a1710 = a1708 & ~l740;
assign a1712 = ~l574 & l572;
assign a1714 = a1712 & a1706;
assign a1716 = a1714 & ~l742;
assign a1718 = ~a1716 & ~a1710;
assign a1720 = ~l578 & ~l576;
assign a1722 = a1720 & a1712;
assign a1724 = a1722 & ~l726;
assign a1726 = l574 & l572;
assign a1728 = a1726 & a1706;
assign a1730 = a1728 & ~i190;
assign a1732 = ~a1730 & ~a1724;
assign a1734 = a1732 & a1718;
assign a1736 = ~l578 & l576;
assign a1738 = a1736 & a1704;
assign a1740 = a1738 & ~l732;
assign a1742 = l574 & ~l572;
assign a1744 = a1742 & a1720;
assign a1746 = a1744 & ~l728;
assign a1748 = ~a1746 & ~a1740;
assign a1750 = l578 & l576;
assign a1752 = a1750 & a1704;
assign a1754 = a1752 & ~i192;
assign a1756 = a1726 & a1720;
assign a1758 = a1756 & ~l730;
assign a1760 = ~a1758 & ~a1754;
assign a1762 = a1760 & a1748;
assign a1764 = a1762 & a1734;
assign a1766 = a1750 & a1726;
assign a1768 = a1766 & ~i188;
assign a1770 = a1750 & a1712;
assign a1772 = a1770 & ~i194;
assign a1774 = ~a1772 & ~a1768;
assign a1776 = a1736 & a1726;
assign a1778 = a1776 & ~l738;
assign a1780 = a1750 & a1742;
assign a1782 = a1780 & ~i196;
assign a1784 = ~a1782 & ~a1778;
assign a1786 = a1784 & a1774;
assign a1788 = a1736 & a1712;
assign a1790 = a1788 & ~l734;
assign a1792 = a1742 & a1706;
assign a1794 = a1792 & ~l744;
assign a1796 = ~a1794 & ~a1790;
assign a1798 = a1742 & a1736;
assign a1800 = a1798 & ~l736;
assign a1802 = a1720 & a1704;
assign a1804 = a1802 & ~l724;
assign a1806 = ~a1804 & ~a1800;
assign a1808 = a1806 & a1796;
assign a1810 = a1808 & a1786;
assign a1812 = a1810 & a1764;
assign a1814 = ~a1812 & l564;
assign a1816 = a1812 & ~l564;
assign a1818 = ~a1816 & ~a1814;
assign a1820 = a1722 & ~l704;
assign a1822 = a1708 & ~l718;
assign a1824 = ~a1822 & ~a1820;
assign a1826 = a1738 & ~l710;
assign a1828 = a1792 & ~l722;
assign a1830 = ~a1828 & ~a1826;
assign a1832 = a1830 & a1824;
assign a1834 = a1728 & ~i180;
assign a1836 = a1798 & ~l714;
assign a1838 = ~a1836 & ~a1834;
assign a1840 = a1788 & ~l712;
assign a1842 = a1770 & ~i184;
assign a1844 = ~a1842 & ~a1840;
assign a1846 = a1844 & a1838;
assign a1848 = a1846 & a1832;
assign a1850 = a1714 & ~l720;
assign a1852 = a1766 & ~i178;
assign a1854 = ~a1852 & ~a1850;
assign a1856 = a1802 & ~l702;
assign a1858 = a1744 & ~l706;
assign a1860 = ~a1858 & ~a1856;
assign a1862 = a1860 & a1854;
assign a1864 = a1752 & ~i182;
assign a1866 = a1780 & ~i186;
assign a1868 = ~a1866 & ~a1864;
assign a1870 = a1756 & ~l708;
assign a1872 = a1776 & ~l716;
assign a1874 = ~a1872 & ~a1870;
assign a1876 = a1874 & a1868;
assign a1878 = a1876 & a1862;
assign a1880 = a1878 & a1848;
assign a1882 = ~a1880 & l562;
assign a1884 = a1880 & ~l562;
assign a1886 = a1798 & ~l692;
assign a1888 = a1738 & ~l688;
assign a1890 = ~a1888 & ~a1886;
assign a1892 = a1788 & ~l690;
assign a1894 = a1752 & ~i172;
assign a1896 = ~a1894 & ~a1892;
assign a1898 = a1896 & a1890;
assign a1900 = a1722 & ~l682;
assign a1902 = a1766 & ~i168;
assign a1904 = ~a1902 & ~a1900;
assign a1906 = a1802 & ~l680;
assign a1908 = a1776 & ~l694;
assign a1910 = ~a1908 & ~a1906;
assign a1912 = a1910 & a1904;
assign a1914 = a1912 & a1898;
assign a1916 = a1728 & ~i170;
assign a1918 = a1714 & ~l698;
assign a1920 = ~a1918 & ~a1916;
assign a1922 = a1792 & ~l700;
assign a1924 = a1708 & ~l696;
assign a1926 = ~a1924 & ~a1922;
assign a1928 = a1926 & a1920;
assign a1930 = a1770 & ~i174;
assign a1932 = a1756 & ~l686;
assign a1934 = ~a1932 & ~a1930;
assign a1936 = a1780 & ~i176;
assign a1938 = a1744 & ~l684;
assign a1940 = ~a1938 & ~a1936;
assign a1942 = a1940 & a1934;
assign a1944 = a1942 & a1928;
assign a1946 = a1944 & a1914;
assign a1948 = ~a1946 & l560;
assign a1950 = a1946 & ~l560;
assign a1952 = a1744 & ~l662;
assign a1954 = a1770 & ~i164;
assign a1956 = ~a1954 & ~a1952;
assign a1958 = a1756 & ~l664;
assign a1960 = a1798 & ~l670;
assign a1962 = ~a1960 & ~a1958;
assign a1964 = a1962 & a1956;
assign a1966 = a1752 & ~i162;
assign a1968 = a1738 & ~l666;
assign a1970 = ~a1968 & ~a1966;
assign a1972 = a1714 & ~l676;
assign a1974 = a1776 & ~l672;
assign a1976 = ~a1974 & ~a1972;
assign a1978 = a1976 & a1970;
assign a1980 = a1978 & a1964;
assign a1982 = a1728 & ~i160;
assign a1984 = a1788 & ~l668;
assign a1986 = ~a1984 & ~a1982;
assign a1988 = a1802 & ~l658;
assign a1990 = a1766 & ~i158;
assign a1992 = ~a1990 & ~a1988;
assign a1994 = a1992 & a1986;
assign a1996 = a1792 & ~l678;
assign a1998 = a1708 & ~l674;
assign a2000 = ~a1998 & ~a1996;
assign a2002 = a1722 & ~l660;
assign a2004 = a1780 & ~i166;
assign a2006 = ~a2004 & ~a2002;
assign a2008 = a2006 & a2000;
assign a2010 = a2008 & a1994;
assign a2012 = a2010 & a1980;
assign a2014 = ~a2012 & l558;
assign a2016 = a2012 & ~l558;
assign a2018 = a1798 & ~l648;
assign a2020 = a1792 & ~l656;
assign a2022 = ~a2020 & ~a2018;
assign a2024 = a1714 & ~l654;
assign a2026 = a1788 & ~l646;
assign a2028 = ~a2026 & ~a2024;
assign a2030 = a2028 & a2022;
assign a2032 = a1756 & ~l642;
assign a2034 = a1708 & ~l652;
assign a2036 = ~a2034 & ~a2032;
assign a2038 = a1802 & ~l636;
assign a2040 = a1744 & ~l640;
assign a2042 = ~a2040 & ~a2038;
assign a2044 = a2042 & a2036;
assign a2046 = a2044 & a2030;
assign a2048 = a1738 & ~l644;
assign a2050 = a1728 & ~i150;
assign a2052 = ~a2050 & ~a2048;
assign a2054 = a1752 & ~i152;
assign a2056 = a1776 & ~l650;
assign a2058 = ~a2056 & ~a2054;
assign a2060 = a2058 & a2052;
assign a2062 = a1766 & ~i148;
assign a2064 = a1722 & ~l638;
assign a2066 = ~a2064 & ~a2062;
assign a2068 = a1770 & ~i154;
assign a2070 = a1780 & ~i156;
assign a2072 = ~a2070 & ~a2068;
assign a2074 = a2072 & a2066;
assign a2076 = a2074 & a2060;
assign a2078 = a2076 & a2046;
assign a2080 = ~a2078 & l556;
assign a2082 = a2078 & ~l556;
assign a2084 = a1708 & ~l632;
assign a2086 = a1738 & ~l624;
assign a2088 = ~a2086 & ~a2084;
assign a2090 = a1752 & ~i142;
assign a2092 = a1792 & ~i138;
assign a2094 = ~a2092 & ~a2090;
assign a2096 = a2094 & a2088;
assign a2098 = a1744 & ~l620;
assign a2100 = a1756 & ~l622;
assign a2102 = ~a2100 & ~a2098;
assign a2104 = a1802 & ~l616;
assign a2106 = a1788 & ~l626;
assign a2108 = ~a2106 & ~a2104;
assign a2110 = a2108 & a2102;
assign a2112 = a2110 & a2096;
assign a2114 = a1776 & ~l630;
assign a2116 = a1766 & ~i136;
assign a2118 = ~a2116 & ~a2114;
assign a2120 = a1728 & ~i140;
assign a2122 = a1770 & ~i144;
assign a2124 = ~a2122 & ~a2120;
assign a2126 = a2124 & a2118;
assign a2128 = a1714 & ~l634;
assign a2130 = a1722 & ~l618;
assign a2132 = ~a2130 & ~a2128;
assign a2134 = a1780 & ~i146;
assign a2136 = a1798 & ~l628;
assign a2138 = ~a2136 & ~a2134;
assign a2140 = a2138 & a2132;
assign a2142 = a2140 & a2126;
assign a2144 = a2142 & a2112;
assign a2146 = ~a2144 & l554;
assign a2148 = a2144 & ~l554;
assign a2150 = a1770 & ~i132;
assign a2152 = a1744 & ~l602;
assign a2154 = ~a2152 & ~a2150;
assign a2156 = a1756 & ~l604;
assign a2158 = a1722 & ~l600;
assign a2160 = ~a2158 & ~a2156;
assign a2162 = a2160 & a2154;
assign a2164 = a1792 & ~i126;
assign a2166 = a1728 & ~i128;
assign a2168 = ~a2166 & ~a2164;
assign a2170 = a1802 & ~l598;
assign a2172 = a1708 & ~l614;
assign a2174 = ~a2172 & ~a2170;
assign a2176 = a2174 & a2168;
assign a2178 = a2176 & a2162;
assign a2180 = a1780 & ~i134;
assign a2182 = a1788 & ~l608;
assign a2184 = ~a2182 & ~a2180;
assign a2186 = a1798 & ~l610;
assign a2188 = a1752 & ~i130;
assign a2190 = ~a2188 & ~a2186;
assign a2192 = a2190 & a2184;
assign a2194 = a1776 & ~l612;
assign a2196 = a1766 & ~i122;
assign a2198 = ~a2196 & ~a2194;
assign a2200 = a1714 & ~i124;
assign a2202 = a1738 & ~l606;
assign a2204 = ~a2202 & ~a2200;
assign a2206 = a2204 & a2198;
assign a2208 = a2206 & a2192;
assign a2210 = a2208 & a2178;
assign a2212 = ~a2210 & l552;
assign a2214 = a2210 & ~l552;
assign a2216 = a1714 & ~i110;
assign a2218 = ~a2216 & ~l550;
assign a2220 = a1738 & ~l594;
assign a2222 = a1788 & ~i104;
assign a2224 = ~a2222 & ~a2220;
assign a2226 = a1798 & ~i106;
assign a2228 = a1728 & ~i114;
assign a2230 = ~a2228 & ~a2226;
assign a2232 = a2230 & a2224;
assign a2234 = a2232 & a2218;
assign a2236 = a1708 & ~i108;
assign a2238 = a1792 & ~i112;
assign a2240 = a1722 & ~l590;
assign a2242 = ~a2240 & ~a2238;
assign a2244 = a2242 & ~a2236;
assign a2246 = a1744 & ~i102;
assign a2248 = a1752 & ~i116;
assign a2250 = ~a2248 & ~a2246;
assign a2252 = a1780 & ~i120;
assign a2254 = a1766 & ~i100;
assign a2256 = ~a2254 & ~a2252;
assign a2258 = a2256 & a2250;
assign a2260 = a1770 & ~i118;
assign a2262 = a1802 & ~l588;
assign a2264 = ~a2262 & ~a2260;
assign a2266 = a1756 & ~l592;
assign a2268 = a1776 & ~l596;
assign a2270 = ~a2268 & ~a2266;
assign a2272 = a2270 & a2264;
assign a2274 = a2272 & a2258;
assign a2276 = a2274 & a2244;
assign a2278 = a2276 & a2234;
assign a2280 = ~a2278 & ~a2214;
assign a2282 = ~a2280 & ~a2212;
assign a2284 = ~a2282 & ~a2148;
assign a2286 = ~a2284 & ~a2146;
assign a2288 = ~a2286 & ~a2082;
assign a2290 = ~a2288 & ~a2080;
assign a2292 = ~a2290 & ~a2016;
assign a2294 = ~a2292 & ~a2014;
assign a2296 = ~a2294 & ~a1950;
assign a2298 = ~a2296 & ~a1948;
assign a2300 = ~a2298 & ~a1884;
assign a2302 = ~a2300 & ~a1882;
assign a2304 = a2302 & ~a1818;
assign a2306 = ~a2302 & a1818;
assign a2308 = ~a2306 & ~a2304;
assign a2310 = a1756 & ~l752;
assign a2312 = a1766 & ~i198;
assign a2314 = ~a2312 & ~a2310;
assign a2316 = a1744 & ~l750;
assign a2318 = a1728 & ~i200;
assign a2320 = ~a2318 & ~a2316;
assign a2322 = a2320 & a2314;
assign a2324 = a1798 & ~l758;
assign a2326 = a1780 & ~i206;
assign a2328 = ~a2326 & ~a2324;
assign a2330 = a1752 & ~i202;
assign a2332 = a1738 & ~l754;
assign a2334 = ~a2332 & ~a2330;
assign a2336 = a2334 & a2328;
assign a2338 = a2336 & a2322;
assign a2340 = a1792 & ~l766;
assign a2342 = a1788 & ~l756;
assign a2344 = ~a2342 & ~a2340;
assign a2346 = a1770 & ~i204;
assign a2348 = a1722 & ~l748;
assign a2350 = ~a2348 & ~a2346;
assign a2352 = a2350 & a2344;
assign a2354 = a1802 & ~l746;
assign a2356 = a1708 & ~l762;
assign a2358 = ~a2356 & ~a2354;
assign a2360 = a1714 & ~l764;
assign a2362 = a1776 & ~l760;
assign a2364 = ~a2362 & ~a2360;
assign a2366 = a2364 & a2358;
assign a2368 = a2366 & a2352;
assign a2370 = a2368 & a2338;
assign a2372 = ~a2370 & l566;
assign a2374 = a2370 & ~l566;
assign a2376 = ~a2374 & ~a2372;
assign a2378 = a2376 & a1816;
assign a2380 = ~a2376 & ~a1816;
assign a2382 = ~a2380 & ~a2378;
assign a2384 = a1728 & ~i210;
assign a2386 = a1780 & ~i216;
assign a2388 = ~a2386 & ~a2384;
assign a2390 = a1792 & ~l788;
assign a2392 = a1714 & ~l786;
assign a2394 = ~a2392 & ~a2390;
assign a2396 = a2394 & a2388;
assign a2398 = a1752 & ~i212;
assign a2400 = a1776 & ~l782;
assign a2402 = ~a2400 & ~a2398;
assign a2404 = a1722 & ~l770;
assign a2406 = a1788 & ~l778;
assign a2408 = ~a2406 & ~a2404;
assign a2410 = a2408 & a2402;
assign a2412 = a2410 & a2396;
assign a2414 = a1744 & ~l772;
assign a2416 = a1802 & ~l768;
assign a2418 = ~a2416 & ~a2414;
assign a2420 = a1770 & ~i214;
assign a2422 = a1798 & ~l780;
assign a2424 = ~a2422 & ~a2420;
assign a2426 = a2424 & a2418;
assign a2428 = a1766 & ~i208;
assign a2430 = a1756 & ~l774;
assign a2432 = ~a2430 & ~a2428;
assign a2434 = a1708 & ~l784;
assign a2436 = a1738 & ~l776;
assign a2438 = ~a2436 & ~a2434;
assign a2440 = a2438 & a2432;
assign a2442 = a2440 & a2426;
assign a2444 = a2442 & a2412;
assign a2446 = ~a2444 & l568;
assign a2448 = a2444 & ~l568;
assign a2450 = ~a2448 & ~a2446;
assign a2452 = a2450 & a2374;
assign a2454 = ~a2450 & ~a2374;
assign a2456 = ~a2454 & ~a2452;
assign a2458 = a2374 & ~a1816;
assign a2460 = ~a2458 & ~a2378;
assign a2462 = a1788 & ~l800;
assign a2464 = a1770 & ~i224;
assign a2466 = ~a2464 & ~a2462;
assign a2468 = a1722 & ~l792;
assign a2470 = a1780 & ~i226;
assign a2472 = ~a2470 & ~a2468;
assign a2474 = a2472 & a2466;
assign a2476 = a1752 & ~i222;
assign a2478 = a1714 & ~l808;
assign a2480 = ~a2478 & ~a2476;
assign a2482 = a1708 & ~l806;
assign a2484 = a1798 & ~l802;
assign a2486 = ~a2484 & ~a2482;
assign a2488 = a2486 & a2480;
assign a2490 = a2488 & a2474;
assign a2492 = a1744 & ~l794;
assign a2494 = a1728 & ~i220;
assign a2496 = ~a2494 & ~a2492;
assign a2498 = a1802 & ~l790;
assign a2500 = a1756 & ~l796;
assign a2502 = ~a2500 & ~a2498;
assign a2504 = a2502 & a2496;
assign a2506 = a1776 & ~l804;
assign a2508 = a1738 & ~l798;
assign a2510 = ~a2508 & ~a2506;
assign a2512 = a1766 & ~i218;
assign a2514 = a1792 & ~l810;
assign a2516 = ~a2514 & ~a2512;
assign a2518 = a2516 & a2510;
assign a2520 = a2518 & a2504;
assign a2522 = a2520 & a2490;
assign a2524 = ~a2522 & l570;
assign a2526 = a2524 & ~a2448;
assign a2528 = ~a2524 & a2448;
assign a2530 = ~a2528 & ~a2526;
assign a2532 = a2522 & ~l570;
assign a2534 = a2448 & ~a2374;
assign a2536 = ~a2534 & ~a2452;
assign a2538 = l816 & l814;
assign a2540 = a2538 & l818;
assign a2542 = a2540 & l820;
assign a2544 = a2542 & l822;
assign a2548 = a2546 & l262;
assign a2550 = l274 & i28;
assign a2552 = ~a2550 & ~a2546;
assign a2554 = a2552 & l246;
assign a2556 = a2554 & ~l838;
assign a2558 = ~a2556 & ~a2548;
assign a2560 = a2546 & l260;
assign a2562 = a2554 & ~l836;
assign a2564 = ~a2562 & ~a2560;
assign a2566 = a2546 & l258;
assign a2568 = a2554 & ~l834;
assign a2570 = ~a2568 & ~a2566;
assign a2572 = a2546 & l256;
assign a2574 = a2554 & l832;
assign a2576 = ~a2574 & ~a2572;
assign a2578 = ~a2552 & ~l254;
assign a2580 = ~a2546 & l254;
assign a2584 = a2582 & ~a2576;
assign a2586 = a2584 & ~a2570;
assign a2588 = a2586 & ~a2564;
assign a2590 = a2588 & ~a2558;
assign a2592 = l274 & i22;
assign a2594 = a2592 & l272;
assign a2596 = l274 & i20;
assign a2598 = ~a2596 & ~a2592;
assign a2600 = a2598 & l250;
assign a2602 = a2600 & ~l844;
assign a2604 = ~a2602 & ~a2594;
assign a2606 = a2592 & l266;
assign a2608 = a2600 & ~l268;
assign a2610 = ~a2608 & ~a2606;
assign a2612 = a2592 & l264;
assign a2614 = a2600 & l840;
assign a2616 = ~a2614 & ~a2612;
assign a2618 = a2598 & ~l252;
assign a2620 = a2592 & l252;
assign a2622 = ~a2620 & ~a2618;
assign a2624 = ~a2622 & ~a2616;
assign a2626 = a2624 & ~a2610;
assign a2628 = a2592 & l270;
assign a2630 = a2600 & ~l842;
assign a2632 = ~a2630 & ~a2628;
assign a2634 = ~a2632 & a2626;
assign a2636 = a2634 & ~a2604;
assign a2638 = ~a2582 & a2576;
assign a2640 = a2546 & l246;
assign a2642 = ~a2640 & ~a2552;
assign a2644 = ~a2642 & a2558;
assign a2646 = a2570 & a2564;
assign a2648 = a2646 & a2644;
assign a2650 = a2648 & a2638;
assign a2652 = ~l370 & ~l364;
assign a2654 = a2652 & l280;
assign a2656 = a1260 & ~l364;
assign a2658 = ~a2656 & ~l416;
assign a2660 = ~l366 & l364;
assign a2662 = ~a2660 & ~a2658;
assign a2664 = a2662 & ~a1266;
assign a2666 = ~a2664 & ~a2654;
assign a2668 = ~a2666 & ~l854;
assign a2670 = ~l852 & ~l850;
assign a2672 = a2670 & a2668;
assign a2674 = ~l848 & ~l846;
assign a2676 = a2674 & a2672;
assign a2678 = l852 & l850;
assign a2680 = a2666 & l854;
assign a2682 = a2680 & a2678;
assign a2684 = ~a2682 & ~a2672;
assign a2686 = a2680 & ~l846;
assign a2688 = ~a2686 & ~a2668;
assign a2690 = a2688 & ~a2684;
assign a2692 = a2592 & ~l248;
assign a2696 = ~a2624 & a2610;
assign a2698 = ~a2696 & ~a2626;
assign a2700 = l428 & l288;
assign a2702 = ~l428 & ~l288;
assign a2706 = ~a2700 & ~l290;
assign a2708 = a2700 & l290;
assign a2714 = l330 & l302;
assign a2716 = a2704 & ~l430;
assign a2718 = a2716 & l290;
assign a2720 = a2718 & ~i76;
assign a2722 = l430 & l288;
assign a2724 = a2722 & ~l290;
assign a2726 = a2724 & ~l320;
assign a2728 = a2722 & l290;
assign a2730 = a2728 & ~i74;
assign a2732 = ~a2730 & ~a2726;
assign a2734 = l430 & ~l288;
assign a2736 = a2734 & ~l290;
assign a2738 = a2736 & ~l324;
assign a2740 = a2734 & l290;
assign a2742 = a2740 & ~i78;
assign a2744 = ~a2742 & ~a2738;
assign a2746 = a2744 & a2732;
assign a2748 = a2746 & ~a2720;
assign a2750 = ~a2704 & ~l430;
assign a2752 = a2750 & a2710;
assign a2754 = a2752 & ~l318;
assign a2756 = a2750 & ~a2710;
assign a2758 = a2756 & ~l326;
assign a2760 = a2716 & ~l290;
assign a2762 = a2760 & ~l322;
assign a2764 = ~a2762 & ~a2758;
assign a2766 = a2764 & ~a2754;
assign a2768 = a2766 & a2748;
assign a2770 = a2768 & a2714;
assign a2772 = ~a2714 & ~l294;
assign a2776 = ~a1022 & ~l998;
assign a2780 = ~a2714 & ~l998;
assign a2782 = a2760 & ~l312;
assign a2784 = a2740 & ~i70;
assign a2786 = a2728 & ~i66;
assign a2788 = ~a2786 & ~a2784;
assign a2790 = a2736 & ~l314;
assign a2792 = a2724 & ~l310;
assign a2794 = ~a2792 & ~a2790;
assign a2796 = a2794 & a2788;
assign a2798 = a2796 & ~a2782;
assign a2800 = a2752 & ~i72;
assign a2802 = a2756 & ~l316;
assign a2804 = a2718 & ~i68;
assign a2806 = ~a2804 & ~a2802;
assign a2808 = a2806 & ~a2800;
assign a2810 = a2808 & a2798;
assign a2812 = ~a2810 & a2714;
assign a2814 = ~a2714 & l300;
assign a2816 = ~a2814 & ~a2812;
assign a2818 = ~a1014 & ~l328;
assign a2820 = ~a2818 & l340;
assign a2822 = ~a2820 & ~l286;
assign a2824 = ~a2822 & ~a1022;
assign a2826 = ~a2824 & ~a2714;
assign a2828 = a2810 & ~a2768;
assign a2830 = a2828 & l330;
assign a2832 = ~a2830 & ~a2826;
assign a2834 = ~a1010 & ~l302;
assign a2836 = a2834 & ~a2824;
assign a2840 = ~l432 & ~l304;
assign a2844 = ~a1026 & l306;
assign a2846 = ~a2844 & ~a1042;
assign a2848 = ~a1028 & l308;
assign a2850 = ~a2848 & ~a1054;
assign a2852 = a1054 & ~l376;
assign a2854 = ~a1054 & l310;
assign a2856 = ~a2854 & ~a2852;
assign a2858 = a1058 & ~l376;
assign a2860 = ~a1058 & l312;
assign a2862 = ~a2860 & ~a2858;
assign a2864 = a1062 & ~l376;
assign a2866 = ~a1062 & l314;
assign a2868 = ~a2866 & ~a2864;
assign a2870 = a1066 & ~l376;
assign a2872 = ~a1066 & l316;
assign a2874 = ~a2872 & ~a2870;
assign a2876 = a1050 & ~l422;
assign a2878 = ~a1050 & l318;
assign a2880 = ~a2878 & ~a2876;
assign a2882 = a1054 & ~l422;
assign a2884 = ~a1054 & l320;
assign a2886 = ~a2884 & ~a2882;
assign a2888 = a1058 & ~l422;
assign a2890 = ~a1058 & l322;
assign a2892 = ~a2890 & ~a2888;
assign a2894 = a1062 & ~l422;
assign a2896 = ~a1062 & l324;
assign a2898 = ~a2896 & ~a2894;
assign a2900 = a1066 & ~l422;
assign a2902 = ~a1066 & l326;
assign a2904 = ~a2902 & ~a2900;
assign a2906 = ~a1018 & ~l340;
assign a2908 = ~a2906 & ~a2770;
assign a2912 = l860 & l826;
assign a2914 = ~a2912 & ~l332;
assign a2918 = l434 & ~l338;
assign a2920 = l274 & i26;
assign a2922 = l274 & i24;
assign a2924 = a2922 & ~a2920;
assign a2926 = a2924 & a2918;
assign a2928 = ~l434 & l338;
assign a2930 = a2928 & ~a2592;
assign a2932 = a2930 & ~l336;
assign a2934 = a2932 & l334;
assign a2936 = ~a2934 & ~a2926;
assign a2938 = ~a2920 & a2918;
assign a2940 = a2938 & ~l334;
assign a2942 = a2940 & l336;
assign a2944 = a2596 & ~a2592;
assign a2946 = a2944 & a2928;
assign a2948 = ~a2946 & ~l1004;
assign a2950 = a2948 & ~a2942;
assign a2952 = a2950 & a2936;
assign a2954 = ~a2928 & ~a2918;
assign a2956 = ~a2954 & a2924;
assign a2958 = a2956 & a2944;
assign a2960 = ~a2922 & ~a2920;
assign a2962 = a2960 & a2598;
assign a2964 = ~a2962 & l1004;
assign a2966 = a2964 & ~a2958;
assign a2968 = ~a2966 & l340;
assign a2970 = a2968 & ~a2952;
assign a2972 = a2944 & ~l436;
assign a2974 = a2972 & l438;
assign a2976 = a2960 & ~l1004;
assign a2978 = l1004 & l434;
assign a2980 = a2978 & a2924;
assign a2982 = ~a2980 & ~a2976;
assign a2984 = ~a2982 & a2974;
assign a2986 = ~a2984 & ~a2970;
assign a2988 = l1004 & l442;
assign a2990 = a2988 & l338;
assign a2992 = a2990 & a2944;
assign a2994 = ~a2924 & l442;
assign a2996 = ~l1004 & l442;
assign a2998 = a2996 & a2598;
assign a3000 = ~a2998 & ~a2994;
assign a3002 = a3000 & ~a2992;
assign a3004 = l434 & l338;
assign a3006 = a3004 & l1004;
assign a3008 = l336 & l334;
assign a3010 = a3008 & a2930;
assign a3012 = ~a3010 & ~a3006;
assign a3014 = a3012 & ~a2946;
assign a3016 = l336 & ~l334;
assign a3018 = a3016 & a3004;
assign a3020 = ~a3018 & ~a2924;
assign a3022 = a3020 & a3014;
assign a3024 = ~a3022 & ~a3002;
assign a3026 = ~a2944 & l440;
assign a3028 = ~l336 & l334;
assign a3030 = a3028 & a3004;
assign a3032 = a3008 & a2938;
assign a3034 = ~a3032 & ~a3006;
assign a3036 = a3034 & ~a2926;
assign a3038 = a3036 & ~a3030;
assign a3040 = ~a3038 & a3026;
assign a3042 = ~a3040 & ~a3024;
assign a3044 = a3042 & a2986;
assign a3046 = a3044 & ~l334;
assign a3048 = ~a2976 & a2974;
assign a3050 = ~l1004 & ~l442;
assign a3052 = ~a3050 & ~a2994;
assign a3054 = a3052 & a2946;
assign a3056 = ~a3054 & ~a3048;
assign a3058 = a3056 & ~a3044;
assign a3062 = a3044 & ~l336;
assign a3064 = a2974 & a2926;
assign a3066 = ~a2964 & ~l442;
assign a3068 = ~a3066 & a3000;
assign a3070 = a2946 & ~l442;
assign a3072 = ~a3070 & ~l440;
assign a3074 = a3072 & a3068;
assign a3076 = ~a3074 & ~a3064;
assign a3078 = a3076 & ~a3044;
assign a3082 = ~a3004 & ~a2932;
assign a3084 = ~a3082 & ~l334;
assign a3086 = ~a3084 & a3014;
assign a3088 = a3086 & ~a2924;
assign a3090 = ~l434 & ~l338;
assign a3092 = ~a3090 & l1004;
assign a3094 = ~a3092 & a2598;
assign a3096 = a3090 & ~l1004;
assign a3098 = a3096 & a2944;
assign a3100 = ~a3098 & a2924;
assign a3102 = a3100 & ~a3094;
assign a3104 = ~a3102 & l442;
assign a3106 = a3104 & ~a3088;
assign a3108 = ~a3004 & ~a2940;
assign a3110 = ~a3108 & ~l336;
assign a3112 = ~a3110 & a3036;
assign a3114 = ~a3112 & a3026;
assign a3116 = l1004 & l340;
assign a3118 = a2924 & a2598;
assign a3120 = a2960 & a2944;
assign a3122 = ~a3120 & ~a3118;
assign a3124 = ~a3122 & a3090;
assign a3126 = ~a3124 & ~a2962;
assign a3128 = ~a3126 & a3116;
assign a3130 = ~a3096 & a2922;
assign a3132 = ~a3092 & ~a2920;
assign a3134 = a3132 & ~a3130;
assign a3136 = a3134 & a2974;
assign a3138 = ~l1004 & l340;
assign a3140 = ~a2946 & ~a2932;
assign a3142 = ~a2940 & ~a2926;
assign a3144 = a3142 & a3140;
assign a3146 = ~a3144 & a3138;
assign a3148 = ~a3146 & ~a3136;
assign a3150 = a3148 & ~a3128;
assign a3152 = a3150 & ~a3114;
assign a3154 = a3152 & ~a3106;
assign a3156 = a3154 & ~l338;
assign a3158 = ~a2928 & ~l1004;
assign a3160 = ~a2944 & a2928;
assign a3162 = ~a3160 & ~a3158;
assign a3164 = a3162 & l336;
assign a3166 = ~a3164 & ~a3000;
assign a3168 = ~a2928 & ~a2924;
assign a3170 = ~a3168 & l336;
assign a3172 = ~a3170 & ~l1004;
assign a3174 = ~a3158 & ~a2944;
assign a3176 = ~a3174 & ~l440;
assign a3178 = a3176 & ~a3172;
assign a3180 = ~a3178 & ~l442;
assign a3182 = ~a3180 & ~a3166;
assign a3184 = ~a2918 & l1004;
assign a3186 = ~a3184 & ~a2926;
assign a3188 = a3026 & l336;
assign a3190 = a3188 & ~a3186;
assign a3192 = a3048 & ~a2924;
assign a3194 = ~a3192 & ~a3190;
assign a3196 = a3194 & ~a3182;
assign a3198 = a3196 & ~a3154;
assign a3202 = a3138 & a3090;
assign a3204 = ~a3202 & ~a3146;
assign a3206 = a3204 & l340;
assign a3208 = a3032 & ~a2922;
assign a3210 = ~a3208 & ~a3006;
assign a3212 = ~a3210 & a3026;
assign a3214 = a3010 & ~a2596;
assign a3216 = ~a3214 & ~a3006;
assign a3218 = ~a3216 & a2994;
assign a3220 = a1496 & l1004;
assign a3222 = a3220 & ~a2924;
assign a3224 = a3222 & ~a2944;
assign a3226 = ~a3224 & ~a3218;
assign a3228 = a3226 & ~a3212;
assign a3230 = a3228 & ~a3206;
assign a3234 = a3232 & ~i52;
assign a3236 = ~a3232 & l344;
assign a3238 = ~a3236 & ~a3234;
assign a3240 = a3232 & ~i64;
assign a3242 = ~a3232 & l346;
assign a3244 = ~a3242 & ~a3240;
assign a3246 = a3232 & ~i4;
assign a3248 = ~a3232 & l348;
assign a3250 = ~a3248 & ~a3246;
assign a3252 = a3232 & i10;
assign a3254 = ~a3232 & l350;
assign a3256 = ~a3254 & ~a3252;
assign a3258 = a3232 & ~i12;
assign a3260 = ~a3232 & l352;
assign a3262 = ~a3260 & ~a3258;
assign a3264 = a3232 & i18;
assign a3266 = ~a3232 & l354;
assign a3268 = ~a3266 & ~a3264;
assign a3270 = a3232 & i2;
assign a3272 = ~a3232 & l356;
assign a3274 = ~a3272 & ~a3270;
assign a3276 = a3232 & i62;
assign a3278 = ~a3232 & l358;
assign a3280 = ~a3278 & ~a3276;
assign a3282 = l418 & l416;
assign a3284 = a3282 & l360;
assign a3286 = ~a3282 & ~l360;
assign a3290 = ~a3284 & l362;
assign a3292 = a3284 & ~l362;
assign a3294 = ~a3292 & ~a3290;
assign a3296 = a1072 & l378;
assign a3298 = a3296 & ~a1240;
assign a3300 = l422 & l376;
assign a3302 = a3300 & l828;
assign a3304 = ~a3302 & l408;
assign a3306 = a3304 & ~a3298;
assign a3308 = a1078 & l422;
assign a3310 = a3308 & a1240;
assign a3312 = ~a3310 & ~l408;
assign a3314 = a1260 & l364;
assign a3316 = a3314 & ~a3312;
assign a3318 = a3316 & ~a3306;
assign a3320 = a1078 & ~l366;
assign a3322 = ~a3320 & ~l364;
assign a3324 = ~a3322 & l368;
assign a3326 = a1324 & a1008;
assign a3328 = ~a2656 & ~a2654;
assign a3330 = a3328 & ~a3326;
assign a3332 = a3330 & ~a3324;
assign a3334 = a3332 & ~a3318;
assign a3336 = a3334 & ~l364;
assign a3338 = a1262 & ~a1238;
assign a3340 = l368 & ~l366;
assign a3342 = a3340 & ~a3308;
assign a3344 = ~a3342 & ~l364;
assign a3346 = a3344 & ~a3338;
assign a3348 = a3314 & ~a3298;
assign a3350 = ~a1070 & l422;
assign a3352 = ~a3350 & l828;
assign a3354 = ~a3352 & ~l370;
assign a3356 = ~a3354 & ~a3348;
assign a3358 = a3356 & ~a3346;
assign a3362 = l828 & l372;
assign a3364 = ~a3362 & a3334;
assign a3366 = a3340 & ~a3310;
assign a3368 = a3340 & l364;
assign a3370 = a1008 & ~l364;
assign a3372 = ~a3370 & ~a3368;
assign a3374 = a3372 & ~l372;
assign a3376 = a3374 & ~a3366;
assign a3378 = a3376 & ~a3364;
assign a3380 = a3364 & ~l366;
assign a3384 = a3364 & ~l368;
assign a3386 = a3340 & a3310;
assign a3388 = a3372 & ~a1260;
assign a3390 = a3388 & ~a3386;
assign a3392 = a3390 & ~a3364;
assign a3396 = ~a3394 & ~a3382;
assign a3400 = a3360 & ~l984;
assign a3404 = ~a3398 & ~a1010;
assign a3406 = a3404 & l376;
assign a3408 = a3398 & ~l986;
assign a3410 = ~a3408 & ~a3406;
assign a3412 = a1078 & l372;
assign a3414 = a3394 & ~a3382;
assign a3416 = a3414 & a3360;
assign a3418 = ~a3416 & l378;
assign a3420 = ~a3418 & ~a3412;
assign a3422 = ~l368 & ~l364;
assign a3424 = ~a3422 & l382;
assign a3426 = ~a3424 & ~a1260;
assign a3430 = a1090 & l424;
assign a3432 = ~a1314 & a1298;
assign a3434 = ~l424 & l388;
assign a3436 = a3434 & ~a3432;
assign a3438 = ~a3436 & ~a3430;
assign a3440 = a1152 & a1084;
assign a3442 = a3440 & ~a1180;
assign a3444 = ~a3440 & ~l392;
assign a3446 = a3444 & ~a1316;
assign a3450 = ~a3414 & ~l394;
assign a3454 = a3382 & ~l394;
assign a3458 = ~a2654 & l398;
assign a3460 = ~a3458 & ~a3412;
assign a3462 = a1228 & a1206;
assign a3464 = a3462 & a1314;
assign a3466 = l392 & l388;
assign a3468 = a3466 & a1142;
assign a3470 = ~a3468 & ~a1102;
assign a3472 = a3470 & ~l396;
assign a3474 = a3472 & ~a3464;
assign a3476 = a3474 & l400;
assign a3478 = ~a3470 & ~l396;
assign a3480 = a3478 & ~l400;
assign a3482 = l398 & l396;
assign a3484 = ~a3482 & ~a3480;
assign a3486 = a3484 & ~a3476;
assign a3488 = a3474 & l402;
assign a3490 = l402 & ~l400;
assign a3492 = ~a3490 & ~a1098;
assign a3494 = a3492 & a3478;
assign a3496 = ~a3494 & ~a3482;
assign a3498 = a3496 & ~a3488;
assign a3500 = ~a3464 & ~a1234;
assign a3502 = ~l402 & ~l382;
assign a3504 = ~a3502 & a1232;
assign a3506 = ~a1316 & ~l406;
assign a3508 = a3506 & ~a3504;
assign a3512 = a3500 & l408;
assign a3514 = a1324 & l406;
assign a3516 = a3514 & a3504;
assign a3518 = ~a3516 & ~a3512;
assign a3520 = ~l420 & l282;
assign a3522 = l422 & ~l408;
assign a3524 = a3522 & ~a3520;
assign a3526 = a1070 & l408;
assign a3528 = ~a3526 & l378;
assign a3530 = a3528 & ~a3524;
assign a3532 = a3530 & ~l410;
assign a3534 = ~a3530 & l410;
assign a3536 = ~a3534 & ~a3532;
assign a3540 = ~a3532 & l412;
assign a3542 = a3532 & ~l412;
assign a3544 = ~a3542 & ~a3540;
assign a3548 = ~a3542 & l414;
assign a3550 = a3532 & a1238;
assign a3552 = ~a3550 & l370;
assign a3554 = a3552 & ~a3548;
assign a3558 = ~l418 & ~l416;
assign a3564 = a3398 & ~l990;
assign a3566 = ~a3564 & ~a3562;
assign a3570 = a3568 & a1170;
assign a3572 = a1316 & ~l278;
assign a3574 = l406 & ~l388;
assign a3576 = a3574 & a1232;
assign a3578 = ~a3576 & ~a3572;
assign a3580 = ~a3578 & l382;
assign a3582 = a3490 & a1092;
assign a3584 = ~a3582 & ~a1144;
assign a3586 = a1148 & a1086;
assign a3588 = a3586 & ~a3584;
assign a3590 = a3582 & l404;
assign a3592 = l390 & l388;
assign a3594 = a3592 & a1098;
assign a3596 = a3594 & a1142;
assign a3598 = ~a3596 & l426;
assign a3600 = a3598 & ~a3590;
assign a3602 = a3600 & ~a3588;
assign a3604 = a3602 & ~a3580;
assign a3606 = ~a3604 & ~a3570;
assign a3610 = ~l430 & ~l302;
assign a3614 = a3352 & a1324;
assign a3616 = ~a3614 & ~l432;
assign a3618 = ~a3616 & a3370;
assign a3620 = a3308 & ~a1238;
assign a3622 = l426 & ~i80;
assign a3624 = a3622 & a3300;
assign a3626 = a3624 & a3314;
assign a3628 = ~a3626 & ~a3620;
assign a3630 = ~a3370 & l406;
assign a3632 = a3630 & ~a3628;
assign a3634 = ~a3632 & ~a3618;
assign a3636 = a3154 & ~l434;
assign a3638 = ~a3186 & l334;
assign a3640 = ~a3638 & l440;
assign a3642 = a3068 & ~a2944;
assign a3644 = ~a3168 & a3050;
assign a3646 = ~a3158 & a2994;
assign a3648 = ~a3646 & ~a3644;
assign a3650 = ~a3648 & ~a3160;
assign a3652 = ~a3650 & ~l440;
assign a3654 = ~a3652 & l334;
assign a3656 = ~a3654 & ~a3642;
assign a3658 = ~a3656 & ~a3640;
assign a3660 = ~a3154 & ~a3048;
assign a3662 = a3660 & ~a3658;
assign a3666 = ~a3104 & ~a2992;
assign a3668 = ~a3090 & a3086;
assign a3670 = a3668 & ~a2924;
assign a3672 = ~a3670 & ~a3666;
assign a3674 = a3112 & ~a3090;
assign a3676 = ~a2944 & ~l436;
assign a3678 = a3676 & ~a3674;
assign a3680 = ~a3134 & ~a2980;
assign a3682 = ~a3680 & a2972;
assign a3684 = ~a3682 & ~a1496;
assign a3686 = a3684 & a3204;
assign a3688 = a3686 & ~a3678;
assign a3690 = a3688 & ~a3672;
assign a3692 = a3116 & a2958;
assign a3694 = ~a3692 & ~a3128;
assign a3696 = a3694 & a3690;
assign a3698 = ~l336 & ~l334;
assign a3700 = ~a3698 & a3160;
assign a3702 = ~l442 & ~l434;
assign a3704 = ~a3702 & a2924;
assign a3706 = l1004 & l438;
assign a3708 = ~a3706 & ~a2978;
assign a3710 = a3708 & ~a3704;
assign a3712 = a3710 & ~a3700;
assign a3714 = a3712 & ~a3696;
assign a3716 = ~a3714 & l436;
assign a3718 = a3698 & a3186;
assign a3720 = ~a3718 & ~a3090;
assign a3722 = ~a3720 & l438;
assign a3724 = ~l1004 & ~l438;
assign a3726 = a3724 & ~a2924;
assign a3728 = ~a3726 & a3676;
assign a3730 = a3728 & ~a3722;
assign a3732 = a3730 & ~a3696;
assign a3734 = ~a3732 & ~a3716;
assign a3736 = a3690 & ~l438;
assign a3738 = ~a3702 & ~a3698;
assign a3740 = ~a3738 & ~a3162;
assign a3742 = ~a3090 & l436;
assign a3744 = a3742 & ~a2924;
assign a3746 = a3744 & ~a3740;
assign a3748 = ~a2948 & l340;
assign a3750 = ~a3748 & ~a2972;
assign a3752 = a3750 & ~a3746;
assign a3754 = a3752 & ~a3696;
assign a3756 = ~a3754 & ~a3736;
assign a3758 = ~a3698 & ~l338;
assign a3760 = a3758 & ~a2924;
assign a3762 = ~a3760 & ~a3184;
assign a3764 = ~a3090 & l440;
assign a3766 = a3764 & ~a3762;
assign a3768 = ~a3766 & ~a3222;
assign a3770 = a3768 & ~a3756;
assign a3772 = ~a3674 & a3026;
assign a3774 = a2942 & ~a2922;
assign a3776 = ~a3774 & ~a2946;
assign a3778 = ~a3776 & a3138;
assign a3780 = a3004 & ~l1004;
assign a3782 = a3780 & a3016;
assign a3784 = ~a3782 & ~a2946;
assign a3786 = ~a3784 & a2994;
assign a3788 = ~a2972 & ~l440;
assign a3790 = a3788 & ~a3786;
assign a3792 = a3790 & ~a3778;
assign a3796 = ~a3668 & ~a2924;
assign a3798 = ~a3796 & l442;
assign a3800 = ~a2926 & a2596;
assign a3802 = ~a3800 & a3138;
assign a3804 = a3802 & ~a2936;
assign a3806 = ~a2944 & a1496;
assign a3808 = a3806 & a2924;
assign a3810 = a3780 & a3028;
assign a3812 = ~a3810 & ~a2926;
assign a3814 = ~a3812 & a3026;
assign a3816 = ~a3814 & ~a3808;
assign a3818 = a3816 & ~a3804;
assign a3820 = a3818 & ~a3798;
assign a3822 = ~a2652 & a1142;
assign a3828 = a3568 & a1142;
assign a3830 = a3490 & a1084;
assign a3832 = a3830 & a1142;
assign a3834 = ~a3832 & l448;
assign a3836 = ~a3834 & ~a3828;
assign a3838 = ~l450 & ~l448;
assign a3840 = ~a3838 & ~a1276;
assign a3844 = ~a1276 & ~l452;
assign a3846 = ~a3844 & ~a1010;
assign a3850 = ~a1278 & ~l454;
assign a3852 = ~a3850 & ~a1010;
assign a3856 = ~a1280 & ~l456;
assign a3858 = ~a3856 & ~a1010;
assign a3862 = ~a1282 & ~l458;
assign a3864 = ~a3862 & ~a1010;
assign a3868 = ~a1284 & ~l460;
assign a3870 = ~a3868 & ~a1010;
assign a3874 = ~a1286 & ~l462;
assign a3876 = ~a3874 & ~a1010;
assign a3880 = ~a1288 & ~l464;
assign a3882 = ~a3880 & ~a1010;
assign a3886 = ~a1290 & ~l466;
assign a3888 = ~a3886 & ~a1010;
assign a3892 = ~a1292 & ~l468;
assign a3894 = ~a3892 & ~a1010;
assign a3898 = ~a1294 & ~l470;
assign a3904 = a1430 & ~a1336;
assign a3906 = ~a3904 & ~a1328;
assign a3908 = a1344 & ~a1332;
assign a3910 = a3908 & ~a3906;
assign a3912 = ~a1372 & l472;
assign a3914 = ~a3912 & a1116;
assign a3916 = ~a1334 & ~l472;
assign a3918 = ~a1344 & ~a1336;
assign a3920 = a3918 & ~a1386;
assign a3922 = a3920 & ~a3916;
assign a3924 = a3922 & ~a3914;
assign a3926 = a3924 & a1428;
assign a3928 = ~a3926 & ~a3910;
assign a3932 = a1118 & l426;
assign a3934 = ~a3902 & l484;
assign a3936 = ~a3934 & ~a3932;
assign a3938 = l274 & i18;
assign a3940 = l274 & i12;
assign a3942 = a3940 & ~a3938;
assign a3944 = l274 & i4;
assign a3946 = a3944 & ~i10;
assign a3948 = ~a3946 & ~a3942;
assign a3950 = l274 & i2;
assign a3952 = l274 & i64;
assign a3954 = ~a3952 & ~a3950;
assign a3956 = l274 & i62;
assign a3958 = l274 & i52;
assign a3960 = ~a3958 & ~a3956;
assign a3962 = ~a3960 & ~a3954;
assign a3964 = a3962 & a3948;
assign a3966 = a3952 & ~a3950;
assign a3968 = ~a3966 & a3948;
assign a3970 = l274 & i10;
assign a3972 = ~a3970 & ~a3944;
assign a3974 = ~a3972 & ~a3942;
assign a3976 = a3974 & ~a3966;
assign a3978 = ~a3976 & ~a3968;
assign a3980 = a3978 & ~a3964;
assign a3984 = ~i92 & i30;
assign a3986 = i94 & ~i34;
assign a3988 = ~a3986 & ~a3984;
assign a3990 = i92 & ~i30;
assign a3992 = ~i94 & i34;
assign a3994 = ~a3992 & ~a3990;
assign a3996 = a3994 & a3988;
assign a3998 = ~a1522 & i96;
assign a4000 = a1522 & ~i96;
assign a4002 = ~a4000 & ~a3998;
assign a4004 = a4002 & a3996;
assign a4006 = a1540 & i98;
assign a4008 = ~a1540 & ~i98;
assign a4010 = ~a4008 & ~a4006;
assign a4012 = ~a4010 & ~a1538;
assign a4014 = a4012 & a4004;
assign a4016 = a4014 & l538;
assign a4018 = a1662 & ~a1552;
assign a4020 = a4018 & ~a4016;
assign a4022 = a3974 & ~a3954;
assign a4024 = a4022 & ~a2552;
assign a4026 = ~a3970 & ~a3950;
assign a4028 = ~a3956 & ~a3938;
assign a4030 = a4028 & a4026;
assign a4032 = ~a4030 & a4022;
assign a4034 = ~a4032 & ~a2546;
assign a4036 = a4034 & i84;
assign a4038 = ~a4036 & i82;
assign a4040 = ~a4038 & a4024;
assign a4042 = a4040 & ~a4020;
assign a4044 = a3938 & ~i4;
assign a4046 = ~a4044 & a4026;
assign a4048 = ~a4046 & a3948;
assign a4050 = ~a4048 & ~a3956;
assign a4052 = a4050 & a3968;
assign a4054 = ~a4030 & a3976;
assign a4056 = ~a4054 & ~a3968;
assign a4058 = ~a4056 & ~a4052;
assign a4060 = ~a4050 & a3964;
assign a4062 = a4060 & a3978;
assign a4064 = ~a4062 & ~a2546;
assign a4066 = a4064 & ~a4058;
assign a4068 = a4066 & i86;
assign a4070 = ~a4068 & l486;
assign a4072 = ~a4070 & a3982;
assign a4074 = ~a4072 & a4042;
assign a4076 = a4072 & a4020;
assign a4078 = ~i90 & ~i88;
assign a4080 = ~a4078 & l490;
assign a4082 = ~a4080 & ~a4040;
assign a4084 = a4082 & a4076;
assign a4086 = ~a4084 & ~a4074;
assign a4088 = ~a4072 & ~a4040;
assign a4090 = ~a4088 & a1538;
assign a4092 = ~a4090 & ~a4086;
assign a4094 = i90 & i88;
assign a4096 = a4094 & ~a4074;
assign a4098 = a4078 & a4074;
assign a4100 = ~a4098 & ~a4096;
assign a4102 = ~a4100 & a4092;
assign a4104 = a4102 & ~l490;
assign a4106 = ~a4102 & l490;
assign a4108 = ~a4106 & ~a4104;
assign a4110 = ~l536 & l512;
assign a4112 = a4110 & a4082;
assign a4114 = a4042 & ~a1624;
assign a4116 = a4114 & a1666;
assign a4118 = ~a4116 & ~a4112;
assign a4120 = a4076 & ~a1538;
assign a4122 = a4120 & ~a4118;
assign a4124 = a4122 & i30;
assign a4126 = ~a4122 & l492;
assign a4128 = ~a4126 & ~a4124;
assign a4130 = a4122 & i34;
assign a4132 = ~a4122 & l494;
assign a4134 = ~a4132 & ~a4130;
assign a4136 = a4122 & a1522;
assign a4138 = ~a4122 & l496;
assign a4140 = ~a4138 & ~a4136;
assign a4142 = a4122 & a1540;
assign a4144 = ~a4122 & l498;
assign a4146 = ~a4144 & ~a4142;
assign a4148 = ~a4110 & ~l500;
assign a4150 = ~a4086 & a1584;
assign a4152 = ~a4150 & l500;
assign a4154 = a4092 & a4076;
assign a4156 = ~a4154 & ~a4152;
assign a4160 = l536 & l512;
assign a4162 = a4160 & a4082;
assign a4164 = a4114 & ~a1666;
assign a4166 = ~a4164 & ~a4162;
assign a4168 = ~a4166 & a4120;
assign a4170 = a4168 & i30;
assign a4172 = ~a4168 & l502;
assign a4174 = ~a4172 & ~a4170;
assign a4176 = a4168 & i34;
assign a4178 = ~a4168 & l504;
assign a4180 = ~a4178 & ~a4176;
assign a4182 = a4168 & a1522;
assign a4184 = ~a4168 & l506;
assign a4186 = ~a4184 & ~a4182;
assign a4188 = a4168 & a1540;
assign a4190 = ~a4168 & l508;
assign a4192 = ~a4190 & ~a4188;
assign a4194 = ~a4086 & a1620;
assign a4196 = ~a4194 & l510;
assign a4198 = ~a4160 & ~l510;
assign a4200 = ~a4198 & a4154;
assign a4202 = ~a4200 & ~a4196;
assign a4204 = ~a4198 & ~a4148;
assign a4206 = l538 & l512;
assign a4208 = a4206 & l534;
assign a4210 = ~a4208 & a4204;
assign a4212 = ~l524 & ~l522;
assign a4214 = ~a4212 & a4154;
assign a4216 = a4214 & ~a4210;
assign a4218 = ~a4092 & l512;
assign a4220 = a4092 & ~a1624;
assign a4222 = ~a4220 & ~a4218;
assign a4224 = a4222 & ~a4216;
assign a4226 = a4042 & a1658;
assign a4228 = a4082 & l524;
assign a4230 = ~a4228 & ~a4226;
assign a4232 = ~a4230 & a4120;
assign a4234 = a4232 & i30;
assign a4236 = ~a4232 & l514;
assign a4238 = ~a4236 & ~a4234;
assign a4240 = a4232 & i34;
assign a4242 = ~a4232 & l516;
assign a4244 = ~a4242 & ~a4240;
assign a4246 = a4232 & a1522;
assign a4248 = ~a4232 & l518;
assign a4250 = ~a4248 & ~a4246;
assign a4252 = a4232 & a1540;
assign a4254 = ~a4232 & l520;
assign a4256 = ~a4254 & ~a4252;
assign a4258 = ~a4086 & a1656;
assign a4260 = ~a4258 & l522;
assign a4262 = ~a4260 & ~a4214;
assign a4264 = ~l524 & ~l512;
assign a4266 = a4264 & ~l536;
assign a4268 = ~a4266 & ~l538;
assign a4270 = ~a4268 & a4076;
assign a4272 = a4264 & l536;
assign a4274 = ~a4272 & ~l534;
assign a4276 = ~a4274 & a4204;
assign a4278 = a4276 & a4270;
assign a4280 = ~a4278 & a4092;
assign a4282 = ~a4280 & l524;
assign a4284 = a4212 & a4076;
assign a4286 = ~a4284 & ~a1658;
assign a4288 = ~a4286 & a4092;
assign a4290 = ~a4288 & ~a4282;
assign a4292 = a4272 & a4082;
assign a4294 = a4040 & a1552;
assign a4296 = ~a4294 & ~a4292;
assign a4298 = ~a4296 & a4120;
assign a4300 = a4298 & i30;
assign a4302 = ~a4298 & l526;
assign a4304 = ~a4302 & ~a4300;
assign a4306 = a4298 & i34;
assign a4308 = ~a4298 & l528;
assign a4310 = ~a4308 & ~a4306;
assign a4312 = a4298 & a1522;
assign a4314 = ~a4298 & l530;
assign a4316 = ~a4314 & ~a4312;
assign a4318 = a4298 & a1540;
assign a4320 = ~a4298 & l532;
assign a4322 = ~a4320 & ~a4318;
assign a4324 = ~a4086 & a1550;
assign a4326 = ~a4324 & l534;
assign a4328 = ~a4326 & ~a4154;
assign a4332 = l538 & l536;
assign a4334 = ~a4332 & ~a4274;
assign a4336 = ~a4334 & ~a4148;
assign a4338 = ~a4336 & ~a4198;
assign a4340 = ~a4338 & a4214;
assign a4342 = ~a4092 & l536;
assign a4344 = a4092 & ~a1666;
assign a4346 = ~a4344 & ~a4342;
assign a4348 = a4346 & ~a4340;
assign a4350 = ~a4086 & a4014;
assign a4352 = ~a4350 & l538;
assign a4354 = a4270 & a4092;
assign a4356 = ~a4354 & ~a4352;
assign a4358 = a2546 & l284;
assign a4360 = ~a2552 & ~l342;
assign a4362 = a4360 & ~a4358;
assign a4364 = ~a4362 & ~l546;
assign a4366 = ~a4364 & a1670;
assign a4368 = a4362 & ~a1678;
assign a4370 = ~a4368 & ~a1670;
assign a4372 = ~a4370 & ~a4366;
assign a4374 = ~a4372 & ~l540;
assign a4376 = a4362 & ~a1670;
assign a4378 = l548 & l540;
assign a4380 = ~a4378 & ~a1672;
assign a4382 = a4380 & a4376;
assign a4384 = ~a4380 & ~a4376;
assign a4386 = ~a4384 & ~a4382;
assign a4388 = ~a4386 & a4372;
assign a4392 = ~a4378 & ~a4376;
assign a4394 = ~a4392 & a4372;
assign a4396 = a4376 & ~a1672;
assign a4398 = ~a4396 & a4394;
assign a4400 = a4398 & ~l542;
assign a4402 = ~a4398 & l542;
assign a4404 = ~a4402 & ~a4400;
assign a4406 = a4376 & ~a1674;
assign a4408 = ~a4376 & ~l542;
assign a4410 = ~a4408 & ~a4406;
assign a4412 = a4410 & a4394;
assign a4414 = ~a4412 & l544;
assign a4416 = a4412 & ~l544;
assign a4418 = ~a4416 & ~a4414;
assign a4420 = ~a4376 & ~l544;
assign a4422 = a4376 & l544;
assign a4424 = ~a4422 & ~a4420;
assign a4426 = a4424 & a4412;
assign a4428 = a4426 & l546;
assign a4430 = ~a4426 & ~l546;
assign a4434 = a4372 & ~l548;
assign a4436 = ~a4372 & l548;
assign a4438 = ~a4436 & ~a4434;
assign a4440 = a1680 & ~l550;
assign a4444 = ~a1682 & ~l552;
assign a4448 = ~a1684 & ~l554;
assign a4452 = ~a1686 & ~l556;
assign a4456 = ~a1688 & ~l558;
assign a4460 = ~a1690 & ~l560;
assign a4464 = ~a1692 & ~l562;
assign a4468 = ~a1694 & ~l564;
assign a4472 = ~a1696 & ~l566;
assign a4476 = ~a1698 & ~l568;
assign a4480 = ~a1700 & ~l570;
assign a4482 = ~a4368 & ~l572;
assign a4484 = a4368 & l572;
assign a4488 = ~a4484 & ~l574;
assign a4490 = a4484 & l574;
assign a4494 = ~a4490 & ~l576;
assign a4496 = a4490 & l576;
assign a4500 = ~a4496 & l578;
assign a4502 = a4368 & a1776;
assign a4504 = ~a4502 & ~a4500;
assign a4506 = ~a4368 & ~a4364;
assign a4508 = ~a4506 & a1670;
assign a4510 = a4508 & l580;
assign a4512 = ~a4508 & ~l580;
assign a4516 = ~a4510 & ~l582;
assign a4518 = a4510 & l582;
assign a4522 = ~a4518 & ~l584;
assign a4524 = a4518 & l584;
assign a4528 = ~l586 & l584;
assign a4530 = a4528 & a4518;
assign a4532 = ~a4524 & l586;
assign a4534 = ~a4532 & ~a4530;
assign a4536 = a4508 & ~l580;
assign a4538 = ~l586 & ~l584;
assign a4540 = a4538 & ~l582;
assign a4542 = a4540 & a4536;
assign a4544 = a4542 & l550;
assign a4546 = ~a4542 & l588;
assign a4548 = ~a4546 & ~a4544;
assign a4550 = a4540 & a4510;
assign a4552 = a4550 & l550;
assign a4554 = ~a4550 & l590;
assign a4556 = ~a4554 & ~a4552;
assign a4558 = a4538 & a4518;
assign a4560 = a4558 & l550;
assign a4562 = ~a4558 & l592;
assign a4564 = ~a4562 & ~a4560;
assign a4566 = a4528 & ~l582;
assign a4568 = a4566 & a4536;
assign a4570 = a4568 & l550;
assign a4572 = ~a4568 & l594;
assign a4574 = ~a4572 & ~a4570;
assign a4576 = a4530 & l550;
assign a4578 = ~a4530 & l596;
assign a4580 = ~a4578 & ~a4576;
assign a4582 = a4542 & l552;
assign a4584 = ~a4542 & l598;
assign a4586 = ~a4584 & ~a4582;
assign a4588 = a4550 & l552;
assign a4590 = ~a4550 & l600;
assign a4592 = ~a4590 & ~a4588;
assign a4594 = a4536 & l582;
assign a4596 = a4594 & a4538;
assign a4598 = a4596 & l552;
assign a4600 = ~a4596 & l602;
assign a4602 = ~a4600 & ~a4598;
assign a4604 = a4558 & l552;
assign a4606 = ~a4558 & l604;
assign a4608 = ~a4606 & ~a4604;
assign a4610 = a4568 & l552;
assign a4612 = ~a4568 & l606;
assign a4614 = ~a4612 & ~a4610;
assign a4616 = a4566 & a4510;
assign a4618 = a4616 & l552;
assign a4620 = ~a4616 & l608;
assign a4622 = ~a4620 & ~a4618;
assign a4624 = a4594 & a4528;
assign a4626 = a4624 & l552;
assign a4628 = ~a4624 & l610;
assign a4630 = ~a4628 & ~a4626;
assign a4632 = a4530 & l552;
assign a4634 = ~a4530 & l612;
assign a4636 = ~a4634 & ~a4632;
assign a4638 = l586 & ~l584;
assign a4640 = a4638 & ~l582;
assign a4642 = a4640 & a4536;
assign a4644 = a4642 & l552;
assign a4646 = ~a4642 & l614;
assign a4648 = ~a4646 & ~a4644;
assign a4650 = a4542 & l554;
assign a4652 = ~a4542 & l616;
assign a4654 = ~a4652 & ~a4650;
assign a4656 = a4550 & l554;
assign a4658 = ~a4550 & l618;
assign a4660 = ~a4658 & ~a4656;
assign a4662 = a4596 & l554;
assign a4664 = ~a4596 & l620;
assign a4666 = ~a4664 & ~a4662;
assign a4668 = a4558 & l554;
assign a4670 = ~a4558 & l622;
assign a4672 = ~a4670 & ~a4668;
assign a4674 = a4568 & l554;
assign a4676 = ~a4568 & l624;
assign a4678 = ~a4676 & ~a4674;
assign a4680 = a4616 & l554;
assign a4682 = ~a4616 & l626;
assign a4684 = ~a4682 & ~a4680;
assign a4686 = a4624 & l554;
assign a4688 = ~a4624 & l628;
assign a4690 = ~a4688 & ~a4686;
assign a4692 = a4530 & l554;
assign a4694 = ~a4530 & l630;
assign a4696 = ~a4694 & ~a4692;
assign a4698 = a4642 & l554;
assign a4700 = ~a4642 & l632;
assign a4702 = ~a4700 & ~a4698;
assign a4704 = a4640 & a4510;
assign a4706 = a4704 & l554;
assign a4708 = ~a4704 & l634;
assign a4710 = ~a4708 & ~a4706;
assign a4712 = a4542 & l556;
assign a4714 = ~a4542 & l636;
assign a4716 = ~a4714 & ~a4712;
assign a4718 = a4550 & l556;
assign a4720 = ~a4550 & l638;
assign a4722 = ~a4720 & ~a4718;
assign a4724 = a4596 & l556;
assign a4726 = ~a4596 & l640;
assign a4728 = ~a4726 & ~a4724;
assign a4730 = a4558 & l556;
assign a4732 = ~a4558 & l642;
assign a4734 = ~a4732 & ~a4730;
assign a4736 = a4568 & l556;
assign a4738 = ~a4568 & l644;
assign a4740 = ~a4738 & ~a4736;
assign a4742 = a4616 & l556;
assign a4744 = ~a4616 & l646;
assign a4746 = ~a4744 & ~a4742;
assign a4748 = a4624 & l556;
assign a4750 = ~a4624 & l648;
assign a4752 = ~a4750 & ~a4748;
assign a4754 = a4530 & l556;
assign a4756 = ~a4530 & l650;
assign a4758 = ~a4756 & ~a4754;
assign a4760 = a4642 & l556;
assign a4762 = ~a4642 & l652;
assign a4764 = ~a4762 & ~a4760;
assign a4766 = a4704 & l556;
assign a4768 = ~a4704 & l654;
assign a4770 = ~a4768 & ~a4766;
assign a4772 = a4638 & a4594;
assign a4774 = a4772 & l556;
assign a4776 = ~a4772 & l656;
assign a4778 = ~a4776 & ~a4774;
assign a4780 = a4542 & l558;
assign a4782 = ~a4542 & l658;
assign a4784 = ~a4782 & ~a4780;
assign a4786 = a4550 & l558;
assign a4788 = ~a4550 & l660;
assign a4790 = ~a4788 & ~a4786;
assign a4792 = a4596 & l558;
assign a4794 = ~a4596 & l662;
assign a4796 = ~a4794 & ~a4792;
assign a4798 = a4558 & l558;
assign a4800 = ~a4558 & l664;
assign a4802 = ~a4800 & ~a4798;
assign a4804 = a4568 & l558;
assign a4806 = ~a4568 & l666;
assign a4808 = ~a4806 & ~a4804;
assign a4810 = a4616 & l558;
assign a4812 = ~a4616 & l668;
assign a4814 = ~a4812 & ~a4810;
assign a4816 = a4624 & l558;
assign a4818 = ~a4624 & l670;
assign a4820 = ~a4818 & ~a4816;
assign a4822 = a4530 & l558;
assign a4824 = ~a4530 & l672;
assign a4826 = ~a4824 & ~a4822;
assign a4828 = a4642 & l558;
assign a4830 = ~a4642 & l674;
assign a4832 = ~a4830 & ~a4828;
assign a4834 = a4704 & l558;
assign a4836 = ~a4704 & l676;
assign a4838 = ~a4836 & ~a4834;
assign a4840 = a4772 & l558;
assign a4842 = ~a4772 & l678;
assign a4844 = ~a4842 & ~a4840;
assign a4846 = a4542 & l560;
assign a4848 = ~a4542 & l680;
assign a4850 = ~a4848 & ~a4846;
assign a4852 = a4550 & l560;
assign a4854 = ~a4550 & l682;
assign a4856 = ~a4854 & ~a4852;
assign a4858 = a4596 & l560;
assign a4860 = ~a4596 & l684;
assign a4862 = ~a4860 & ~a4858;
assign a4864 = a4558 & l560;
assign a4866 = ~a4558 & l686;
assign a4868 = ~a4866 & ~a4864;
assign a4870 = a4568 & l560;
assign a4872 = ~a4568 & l688;
assign a4874 = ~a4872 & ~a4870;
assign a4876 = a4616 & l560;
assign a4878 = ~a4616 & l690;
assign a4880 = ~a4878 & ~a4876;
assign a4882 = a4624 & l560;
assign a4884 = ~a4624 & l692;
assign a4886 = ~a4884 & ~a4882;
assign a4888 = a4530 & l560;
assign a4890 = ~a4530 & l694;
assign a4892 = ~a4890 & ~a4888;
assign a4894 = a4642 & l560;
assign a4896 = ~a4642 & l696;
assign a4898 = ~a4896 & ~a4894;
assign a4900 = a4704 & l560;
assign a4902 = ~a4704 & l698;
assign a4904 = ~a4902 & ~a4900;
assign a4906 = a4772 & l560;
assign a4908 = ~a4772 & l700;
assign a4910 = ~a4908 & ~a4906;
assign a4912 = a4542 & l562;
assign a4914 = ~a4542 & l702;
assign a4916 = ~a4914 & ~a4912;
assign a4918 = a4550 & l562;
assign a4920 = ~a4550 & l704;
assign a4922 = ~a4920 & ~a4918;
assign a4924 = a4596 & l562;
assign a4926 = ~a4596 & l706;
assign a4928 = ~a4926 & ~a4924;
assign a4930 = a4558 & l562;
assign a4932 = ~a4558 & l708;
assign a4934 = ~a4932 & ~a4930;
assign a4936 = a4568 & l562;
assign a4938 = ~a4568 & l710;
assign a4940 = ~a4938 & ~a4936;
assign a4942 = a4616 & l562;
assign a4944 = ~a4616 & l712;
assign a4946 = ~a4944 & ~a4942;
assign a4948 = a4624 & l562;
assign a4950 = ~a4624 & l714;
assign a4952 = ~a4950 & ~a4948;
assign a4954 = a4530 & l562;
assign a4956 = ~a4530 & l716;
assign a4958 = ~a4956 & ~a4954;
assign a4960 = a4642 & l562;
assign a4962 = ~a4642 & l718;
assign a4964 = ~a4962 & ~a4960;
assign a4966 = a4704 & l562;
assign a4968 = ~a4704 & l720;
assign a4970 = ~a4968 & ~a4966;
assign a4972 = a4772 & l562;
assign a4974 = ~a4772 & l722;
assign a4976 = ~a4974 & ~a4972;
assign a4978 = a4542 & l564;
assign a4980 = ~a4542 & l724;
assign a4982 = ~a4980 & ~a4978;
assign a4984 = a4550 & l564;
assign a4986 = ~a4550 & l726;
assign a4988 = ~a4986 & ~a4984;
assign a4990 = a4596 & l564;
assign a4992 = ~a4596 & l728;
assign a4994 = ~a4992 & ~a4990;
assign a4996 = a4558 & l564;
assign a4998 = ~a4558 & l730;
assign a5000 = ~a4998 & ~a4996;
assign a5002 = a4568 & l564;
assign a5004 = ~a4568 & l732;
assign a5006 = ~a5004 & ~a5002;
assign a5008 = a4616 & l564;
assign a5010 = ~a4616 & l734;
assign a5012 = ~a5010 & ~a5008;
assign a5014 = a4624 & l564;
assign a5016 = ~a4624 & l736;
assign a5018 = ~a5016 & ~a5014;
assign a5020 = a4530 & l564;
assign a5022 = ~a4530 & l738;
assign a5024 = ~a5022 & ~a5020;
assign a5026 = a4642 & l564;
assign a5028 = ~a4642 & l740;
assign a5030 = ~a5028 & ~a5026;
assign a5032 = a4704 & l564;
assign a5034 = ~a4704 & l742;
assign a5036 = ~a5034 & ~a5032;
assign a5038 = a4772 & l564;
assign a5040 = ~a4772 & l744;
assign a5042 = ~a5040 & ~a5038;
assign a5044 = a4542 & l566;
assign a5046 = ~a4542 & l746;
assign a5048 = ~a5046 & ~a5044;
assign a5050 = a4550 & l566;
assign a5052 = ~a4550 & l748;
assign a5054 = ~a5052 & ~a5050;
assign a5056 = a4596 & l566;
assign a5058 = ~a4596 & l750;
assign a5060 = ~a5058 & ~a5056;
assign a5062 = a4558 & l566;
assign a5064 = ~a4558 & l752;
assign a5066 = ~a5064 & ~a5062;
assign a5068 = a4568 & l566;
assign a5070 = ~a4568 & l754;
assign a5072 = ~a5070 & ~a5068;
assign a5074 = a4616 & l566;
assign a5076 = ~a4616 & l756;
assign a5078 = ~a5076 & ~a5074;
assign a5080 = a4624 & l566;
assign a5082 = ~a4624 & l758;
assign a5084 = ~a5082 & ~a5080;
assign a5086 = a4530 & l566;
assign a5088 = ~a4530 & l760;
assign a5090 = ~a5088 & ~a5086;
assign a5092 = a4642 & l566;
assign a5094 = ~a4642 & l762;
assign a5096 = ~a5094 & ~a5092;
assign a5098 = a4704 & l566;
assign a5100 = ~a4704 & l764;
assign a5102 = ~a5100 & ~a5098;
assign a5104 = a4772 & l566;
assign a5106 = ~a4772 & l766;
assign a5108 = ~a5106 & ~a5104;
assign a5110 = a4542 & l568;
assign a5112 = ~a4542 & l768;
assign a5114 = ~a5112 & ~a5110;
assign a5116 = a4550 & l568;
assign a5118 = ~a4550 & l770;
assign a5120 = ~a5118 & ~a5116;
assign a5122 = a4596 & l568;
assign a5124 = ~a4596 & l772;
assign a5126 = ~a5124 & ~a5122;
assign a5128 = a4558 & l568;
assign a5130 = ~a4558 & l774;
assign a5132 = ~a5130 & ~a5128;
assign a5134 = a4568 & l568;
assign a5136 = ~a4568 & l776;
assign a5138 = ~a5136 & ~a5134;
assign a5140 = a4616 & l568;
assign a5142 = ~a4616 & l778;
assign a5144 = ~a5142 & ~a5140;
assign a5146 = a4624 & l568;
assign a5148 = ~a4624 & l780;
assign a5150 = ~a5148 & ~a5146;
assign a5152 = a4530 & l568;
assign a5154 = ~a4530 & l782;
assign a5156 = ~a5154 & ~a5152;
assign a5158 = a4642 & l568;
assign a5160 = ~a4642 & l784;
assign a5162 = ~a5160 & ~a5158;
assign a5164 = a4704 & l568;
assign a5166 = ~a4704 & l786;
assign a5168 = ~a5166 & ~a5164;
assign a5170 = a4772 & l568;
assign a5172 = ~a4772 & l788;
assign a5174 = ~a5172 & ~a5170;
assign a5176 = a4542 & l570;
assign a5178 = ~a4542 & l790;
assign a5180 = ~a5178 & ~a5176;
assign a5182 = a4550 & l570;
assign a5184 = ~a4550 & l792;
assign a5186 = ~a5184 & ~a5182;
assign a5188 = a4596 & l570;
assign a5190 = ~a4596 & l794;
assign a5192 = ~a5190 & ~a5188;
assign a5194 = a4558 & l570;
assign a5196 = ~a4558 & l796;
assign a5198 = ~a5196 & ~a5194;
assign a5200 = a4568 & l570;
assign a5202 = ~a4568 & l798;
assign a5204 = ~a5202 & ~a5200;
assign a5206 = a4616 & l570;
assign a5208 = ~a4616 & l800;
assign a5210 = ~a5208 & ~a5206;
assign a5212 = a4624 & l570;
assign a5214 = ~a4624 & l802;
assign a5216 = ~a5214 & ~a5212;
assign a5218 = a4530 & l570;
assign a5220 = ~a4530 & l804;
assign a5222 = ~a5220 & ~a5218;
assign a5224 = a4642 & l570;
assign a5226 = ~a4642 & l806;
assign a5228 = ~a5226 & ~a5224;
assign a5230 = a4704 & l570;
assign a5232 = ~a4704 & l808;
assign a5234 = ~a5232 & ~a5230;
assign a5236 = a4772 & l570;
assign a5238 = ~a4772 & l810;
assign a5240 = ~a5238 & ~a5236;
assign a5242 = a2944 & ~l248;
assign a5244 = ~a5242 & ~l812;
assign a5246 = ~a2944 & ~l814;
assign a5248 = ~a2592 & l814;
assign a5252 = a2592 & l816;
assign a5254 = a2944 & l248;
assign a5256 = ~l816 & ~l814;
assign a5258 = ~a5256 & ~a2538;
assign a5260 = a5258 & a5254;
assign a5262 = ~a5260 & ~a5252;
assign a5264 = ~a2538 & ~l818;
assign a5266 = ~a5264 & ~a2540;
assign a5268 = ~a5266 & l812;
assign a5270 = ~a5268 & a5254;
assign a5272 = a2592 & l818;
assign a5274 = ~a5272 & ~a5270;
assign a5276 = ~a2540 & ~l820;
assign a5278 = ~a5276 & ~a2542;
assign a5280 = ~a5278 & l812;
assign a5282 = ~a5280 & a5254;
assign a5284 = a2592 & l820;
assign a5286 = ~a5284 & ~a5282;
assign a5288 = a2592 & l822;
assign a5290 = ~a5288 & ~a5254;
assign a5292 = ~l822 & l812;
assign a5294 = a5292 & ~a2542;
assign a5302 = ~l992 & ~l982;
assign a5304 = a5302 & ~l988;
assign a5306 = a5304 & a3400;
assign a5308 = ~a5306 & a3396;
assign a5314 = ~a2584 & a2570;
assign a5316 = ~a5314 & ~a2586;
assign a5318 = ~a2586 & a2564;
assign a5320 = ~a5318 & ~a2588;
assign a5324 = a2622 & a2616;
assign a5328 = a2632 & ~a2626;
assign a5330 = ~a5328 & ~a2634;
assign a5334 = ~a2682 & ~l846;
assign a5336 = a2672 & ~l848;
assign a5338 = ~a5336 & ~a2674;
assign a5342 = ~a2684 & l848;
assign a5344 = a2684 & ~l848;
assign a5348 = ~a2688 & l850;
assign a5350 = a2688 & ~l850;
assign a5354 = ~a2678 & ~a2670;
assign a5356 = ~a5350 & ~a2686;
assign a5358 = a5356 & a5354;
assign a5360 = ~a5356 & ~a5354;
assign a5364 = l274 & i16;
assign a5366 = ~a5364 & i14;
assign a5368 = ~a3944 & ~l854;
assign a5370 = a5368 & ~a3940;
assign a5372 = a5370 & a5366;
assign a5374 = a5372 & a4030;
assign a5376 = a5374 & a3240;
assign a5378 = ~a5376 & ~l980;
assign a5380 = a3952 & a3234;
assign a5382 = a5380 & a5374;
assign a5384 = ~l978 & ~l856;
assign a5386 = a5384 & ~a5382;
assign a5388 = ~a4052 & a3958;
assign a5390 = a5366 & a3232;
assign a5392 = a4030 & a3976;
assign a5394 = ~a5392 & ~a3958;
assign a5396 = ~a5394 & a5390;
assign a5398 = a5396 & ~a5388;
assign a5400 = ~a5398 & ~l854;
assign a5402 = ~a5400 & a5386;
assign a5404 = a5390 & a3958;
assign a5406 = a5404 & a5392;
assign a5408 = ~a5406 & ~l854;
assign a5410 = ~a5408 & a5386;
assign a5412 = ~a5410 & ~a5402;
assign a5414 = a5412 & a5378;
assign a5416 = a5402 & a5378;
assign a5418 = ~a5416 & ~a5412;
assign a5420 = a5416 & ~a5408;
assign a5422 = ~a5420 & ~a5414;
assign a5426 = a5422 & ~a2912;
assign a5428 = a2670 & ~l856;
assign a5430 = a5428 & a2674;
assign a5432 = a5430 & a5414;
assign a5434 = ~a5432 & ~a5426;
assign a5436 = ~l860 & ~l826;
assign a5438 = a5436 & l858;
assign a5440 = a5438 & a5422;
assign a5442 = ~a5440 & ~a5434;
assign a5446 = l862 & l854;
assign a5448 = ~l862 & ~l854;
assign a5452 = a5446 & ~l864;
assign a5454 = ~a5446 & l864;
assign a5456 = ~a5454 & ~a5452;
assign a5458 = a5446 & l864;
assign a5460 = a5458 & l866;
assign a5462 = ~a5458 & ~l866;
assign a5466 = l854 & l358;
assign a5468 = ~a5466 & a5460;
assign a5470 = ~a5460 & ~l868;
assign a5474 = a5452 & l866;
assign a5476 = a5474 & ~a5466;
assign a5478 = ~a5474 & ~l870;
assign a5482 = ~l862 & l854;
assign a5484 = a5482 & ~l864;
assign a5486 = a5484 & l866;
assign a5488 = a5486 & ~a5466;
assign a5490 = ~a5486 & ~l872;
assign a5494 = a5458 & ~l866;
assign a5496 = a5494 & ~a5466;
assign a5498 = ~a5494 & ~l874;
assign a5502 = a5482 & l864;
assign a5504 = a5502 & ~l866;
assign a5506 = a5504 & ~a5466;
assign a5508 = ~a5504 & ~l876;
assign a5512 = a5452 & ~l866;
assign a5514 = a5512 & ~a5466;
assign a5516 = ~a5512 & ~l878;
assign a5520 = a5484 & ~l866;
assign a5522 = a5520 & ~a5466;
assign a5524 = ~a5520 & ~l880;
assign a5528 = l854 & ~l346;
assign a5530 = ~a5528 & a5460;
assign a5532 = ~a5460 & ~l882;
assign a5536 = ~a5528 & a5474;
assign a5538 = ~a5474 & ~l884;
assign a5542 = ~a5528 & a5486;
assign a5544 = ~a5486 & ~l886;
assign a5548 = ~a5528 & a5494;
assign a5550 = ~a5494 & ~l888;
assign a5554 = ~a5528 & a5504;
assign a5556 = ~a5504 & ~l890;
assign a5560 = ~a5528 & a5512;
assign a5562 = ~a5512 & ~l892;
assign a5566 = ~a5528 & a5520;
assign a5568 = ~a5520 & ~l894;
assign a5572 = l854 & l356;
assign a5574 = ~a5572 & a5460;
assign a5576 = ~a5460 & ~l896;
assign a5580 = ~a5572 & a5474;
assign a5582 = ~a5474 & ~l898;
assign a5586 = ~a5572 & a5486;
assign a5588 = ~a5486 & ~l900;
assign a5592 = ~a5572 & a5494;
assign a5594 = ~a5494 & ~l902;
assign a5598 = ~a5572 & a5504;
assign a5600 = ~a5504 & ~l904;
assign a5604 = ~a5572 & a5512;
assign a5606 = ~a5512 & ~l906;
assign a5610 = ~a5572 & a5520;
assign a5612 = ~a5520 & ~l908;
assign a5616 = l854 & ~l348;
assign a5618 = ~a5616 & a5474;
assign a5620 = ~a5474 & ~l910;
assign a5624 = ~a5616 & a5486;
assign a5626 = ~a5486 & ~l912;
assign a5630 = ~a5616 & a5494;
assign a5632 = ~a5494 & ~l914;
assign a5636 = ~a5616 & a5504;
assign a5638 = ~a5504 & ~l916;
assign a5642 = ~a5616 & a5512;
assign a5644 = ~a5512 & ~l918;
assign a5648 = ~a5616 & a5520;
assign a5650 = ~a5520 & ~l920;
assign a5654 = l854 & l350;
assign a5656 = ~a5654 & a5460;
assign a5658 = ~a5460 & ~l922;
assign a5662 = ~a5654 & a5474;
assign a5664 = ~a5474 & ~l924;
assign a5668 = ~a5654 & a5486;
assign a5670 = ~a5486 & ~l926;
assign a5674 = ~a5654 & a5494;
assign a5676 = ~a5494 & ~l928;
assign a5680 = ~a5654 & a5504;
assign a5682 = ~a5504 & ~l930;
assign a5686 = ~a5654 & a5512;
assign a5688 = ~a5512 & ~l932;
assign a5692 = ~a5654 & a5520;
assign a5694 = ~a5520 & ~l934;
assign a5698 = l854 & l354;
assign a5700 = ~a5698 & a5460;
assign a5702 = ~a5460 & ~l936;
assign a5706 = ~a5698 & a5474;
assign a5708 = ~a5474 & ~l938;
assign a5712 = ~a5698 & a5486;
assign a5714 = ~a5486 & ~l940;
assign a5718 = ~a5698 & a5494;
assign a5720 = ~a5494 & ~l942;
assign a5724 = ~a5698 & a5504;
assign a5726 = ~a5504 & ~l944;
assign a5730 = ~a5698 & a5512;
assign a5732 = ~a5512 & ~l946;
assign a5736 = ~a5698 & a5520;
assign a5738 = ~a5520 & ~l948;
assign a5742 = l854 & ~l352;
assign a5744 = ~a5742 & a5460;
assign a5746 = ~a5460 & ~l950;
assign a5750 = ~a5742 & a5474;
assign a5752 = ~a5474 & ~l952;
assign a5756 = ~a5742 & a5486;
assign a5758 = ~a5486 & ~l954;
assign a5762 = ~a5742 & a5494;
assign a5764 = ~a5494 & ~l956;
assign a5768 = ~a5742 & a5504;
assign a5770 = ~a5504 & ~l958;
assign a5774 = ~a5742 & a5512;
assign a5776 = ~a5512 & ~l960;
assign a5780 = ~a5742 & a5520;
assign a5782 = ~a5520 & ~l962;
assign a5786 = l854 & ~l344;
assign a5788 = ~a5786 & a5460;
assign a5790 = ~a5460 & ~l964;
assign a5794 = ~a5786 & a5474;
assign a5796 = ~a5474 & ~l966;
assign a5800 = ~a5786 & a5486;
assign a5802 = ~a5486 & ~l968;
assign a5806 = ~a5786 & a5494;
assign a5808 = ~a5494 & ~l970;
assign a5812 = ~a5786 & a5504;
assign a5814 = ~a5504 & ~l972;
assign a5818 = ~a5786 & a5512;
assign a5820 = ~a5512 & ~l974;
assign a5824 = ~a5786 & a5520;
assign a5826 = ~a5520 & ~l976;
assign a5830 = ~a5416 & ~a2912;
assign a5832 = a5410 & ~a2916;
assign a5836 = ~a3560 & a3288;
assign a5838 = a5836 & ~l362;
assign a5840 = a5838 & ~l876;
assign a5842 = a5836 & l362;
assign a5844 = a5842 & ~i228;
assign a5846 = ~a5844 & ~a5840;
assign a5848 = ~a3560 & ~a3288;
assign a5850 = a5848 & ~a3294;
assign a5852 = a5850 & ~l872;
assign a5854 = a3560 & ~a3288;
assign a5856 = a5854 & a3294;
assign a5858 = a5856 & ~l878;
assign a5860 = ~a5858 & ~a5852;
assign a5862 = a5860 & a5846;
assign a5864 = a5854 & ~a3294;
assign a5866 = a5864 & ~l870;
assign a5868 = a3560 & a3288;
assign a5870 = a5868 & l362;
assign a5872 = a5870 & ~l868;
assign a5874 = ~a5872 & ~a5866;
assign a5876 = a5848 & a3294;
assign a5878 = a5876 & ~l880;
assign a5880 = a5868 & ~l362;
assign a5882 = a5880 & ~l874;
assign a5884 = ~a5882 & ~a5878;
assign a5886 = a5884 & a5874;
assign a5890 = a5838 & ~l890;
assign a5892 = a5864 & ~l884;
assign a5894 = ~a5892 & ~a5890;
assign a5896 = a5856 & ~l892;
assign a5898 = a5850 & ~l886;
assign a5900 = ~a5898 & ~a5896;
assign a5902 = a5900 & a5894;
assign a5904 = a5876 & ~l894;
assign a5906 = a5870 & ~l882;
assign a5908 = ~a5906 & ~a5904;
assign a5910 = a5842 & ~i230;
assign a5912 = a5880 & ~l888;
assign a5914 = ~a5912 & ~a5910;
assign a5916 = a5914 & a5908;
assign a5920 = a5870 & ~i234;
assign a5922 = a5842 & ~i236;
assign a5924 = ~a5922 & ~a5920;
assign a5926 = a5856 & ~l918;
assign a5928 = a5838 & ~l916;
assign a5930 = ~a5928 & ~a5926;
assign a5932 = a5930 & a5924;
assign a5934 = a5880 & ~l914;
assign a5936 = a5850 & ~l912;
assign a5938 = ~a5936 & ~a5934;
assign a5940 = a5876 & ~l920;
assign a5942 = a5864 & ~l910;
assign a5944 = ~a5942 & ~a5940;
assign a5946 = a5944 & a5938;
assign a5950 = a5870 & ~l922;
assign a5952 = a5850 & ~l926;
assign a5954 = ~a5952 & ~a5950;
assign a5956 = a5864 & ~l924;
assign a5958 = a5838 & ~l930;
assign a5960 = ~a5958 & ~a5956;
assign a5962 = a5960 & a5954;
assign a5964 = a5856 & ~l932;
assign a5966 = a5876 & ~l934;
assign a5968 = ~a5966 & ~a5964;
assign a5970 = a5842 & ~i238;
assign a5972 = a5880 & ~l928;
assign a5974 = ~a5972 & ~a5970;
assign a5976 = a5974 & a5968;
assign a5980 = a5880 & ~l970;
assign a5982 = a5870 & ~l964;
assign a5984 = ~a5982 & ~a5980;
assign a5986 = a5850 & ~l968;
assign a5988 = a5842 & ~i244;
assign a5990 = ~a5988 & ~a5986;
assign a5992 = a5990 & a5984;
assign a5994 = a5856 & ~l974;
assign a5996 = a5864 & ~l966;
assign a5998 = ~a5996 & ~a5994;
assign a6000 = a5838 & ~l972;
assign a6002 = a5876 & ~l976;
assign a6004 = ~a6002 & ~a6000;
assign a6006 = a6004 & a5998;
assign a6010 = a5870 & ~l896;
assign a6012 = a5876 & ~l908;
assign a6014 = ~a6012 & ~a6010;
assign a6016 = a5880 & ~l902;
assign a6018 = a5842 & ~i232;
assign a6020 = ~a6018 & ~a6016;
assign a6022 = a6020 & a6014;
assign a6024 = a5864 & ~l898;
assign a6026 = a5838 & ~l904;
assign a6028 = ~a6026 & ~a6024;
assign a6030 = a5850 & ~l900;
assign a6032 = a5856 & ~l906;
assign a6034 = ~a6032 & ~a6030;
assign a6036 = a6034 & a6028;
assign a6038 = a6036 & a6022;
assign a6040 = a5850 & ~l954;
assign a6042 = a5870 & ~l950;
assign a6044 = ~a6042 & ~a6040;
assign a6046 = a5842 & ~i242;
assign a6048 = a5838 & ~l958;
assign a6050 = ~a6048 & ~a6046;
assign a6052 = a6050 & a6044;
assign a6054 = a5864 & ~l952;
assign a6056 = a5876 & ~l962;
assign a6058 = ~a6056 & ~a6054;
assign a6060 = a5880 & ~l956;
assign a6062 = a5856 & ~l960;
assign a6064 = ~a6062 & ~a6060;
assign a6066 = a6064 & a6058;
assign a6068 = a6066 & a6052;
assign a6070 = a5880 & ~l942;
assign a6072 = a5876 & ~l948;
assign a6074 = ~a6072 & ~a6070;
assign a6076 = a5856 & ~l946;
assign a6078 = a5838 & ~l944;
assign a6080 = ~a6078 & ~a6076;
assign a6082 = a6080 & a6074;
assign a6084 = a5850 & ~l940;
assign a6086 = a5864 & ~l938;
assign a6088 = ~a6086 & ~a6084;
assign a6090 = a5870 & ~l936;
assign a6092 = a5842 & ~i240;
assign a6094 = ~a6092 & ~a6090;
assign a6096 = a6094 & a6088;
assign a6098 = a6096 & a6082;
assign a6100 = ~a6098 & ~a6068;
assign a6102 = a6100 & ~a6038;
assign a6104 = ~a3230 & ~l340;
assign a6108 = a2908 & ~a2780;
assign a6118 = ~l328 & ~l298;
assign a6120 = ~a2820 & ~l292;
assign a6122 = ~a6120 & ~a1022;
assign a6124 = ~a6122 & ~a6118;
assign a6126 = a6124 & l1004;
assign a6128 = l328 & l298;
assign a6130 = ~a2828 & a2714;
assign a6132 = ~a6130 & ~a6128;
assign a6134 = a6132 & ~a6116;
assign a6136 = ~a6134 & ~a6124;
assign a6138 = ~a6136 & ~a6126;
assign a6140 = ~a6104 & l1006;
assign a6142 = ~a6122 & ~l330;
assign a6144 = ~a6142 & ~l1004;
assign a6146 = a6144 & ~a6134;
assign a6148 = ~a6146 & ~a6140;
assign p0 = c0;
assign c0 = 0;
assign p1 = c0;
assign p2 = c0;
assign p3 = c0;
assign p4 = c0;
assign p5 = c0;
assign p6 = c0;
assign p7 = c0;
assign p8 = c0;
assign p9 = c0;
assign p10 = c0;
assign p11 = c0;
assign p12 = c0;
assign p13 = c0;
assign p14 = c0;
assign p15 = c0;
assign p16 = c0;
assign p17 = c0;
assign p18 = c0;
assign p19 = c0;
assign p20 = c0;
assign p21 = c0;
assign p22 = c0;
assign p23 = c0;
assign p24 = c0;
assign p25 = c0;
assign p26 = c0;
assign p27 = c0;
assign p28 = c0;
assign p29 = c0;
assign p30 = c0;
assign p31 = c0;
assign p32 = c0;
assign p33 = c0;
assign p34 = c0;
assign p35 = c0;
assign p36 = c0;
assign p37 = c0;
assign p38 = c0;
assign p39 = c0;
assign p40 = c0;
assign p41 = c0;
assign p42 = c0;
assign p43 = c0;
assign p44 = c0;
assign p45 = c0;
assign p46 = c0;
assign p47 = c0;
assign p48 = c0;
assign p49 = c0;
assign p50 = c0;
assign p51 = c0;
assign p52 = c0;
assign p53 = c0;
assign p54 = c0;
assign p55 = c0;
assign p56 = c0;
assign p57 = c0;
assign p58 = c0;
assign p59 = c0;
assign p60 = c0;
assign p61 = c0;
assign p62 = c0;
assign p63 = c0;
assign p64 = c0;
assign p65 = c0;
assign p66 = c0;
assign p67 = c0;
assign p68 = c0;
assign p69 = c0;
assign p70 = c0;
assign p71 = c0;
assign p72 = c0;
assign p73 = c0;
assign p74 = c0;
assign p75 = c0;
assign p76 = c0;
assign p77 = c0;
assign p78 = c0;
assign p79 = c0;
assign p80 = c0;
assign p81 = c0;
assign p82 = c0;
assign p83 = c0;
assign p84 = c0;
assign p85 = c0;
assign p86 = c0;
assign p87 = c0;
assign p88 = c0;
assign p89 = c0;
assign p90 = c0;
assign p91 = c0;
assign p92 = c0;
assign p93 = c0;
assign p94 = c0;
assign p95 = c0;
assign p96 = c0;
assign p97 = c0;
assign p98 = c0;
assign p99 = c0;
assign p100 = c0;
assign p101 = c0;
assign p102 = c0;
assign p103 = c0;
assign p104 = c0;
assign p105 = c0;
assign p106 = c0;
assign p107 = c0;
assign p108 = c0;
assign p109 = c0;
assign p110 = c0;
assign p111 = c0;
assign p112 = c0;
assign p113 = c0;
assign p114 = c0;
assign p115 = c0;
assign p116 = c0;
assign p117 = c0;
assign p118 = c0;
assign p119 = c0;
assign p120 = c0;
assign p121 = c0;
assign p122 = c0;
assign p123 = c0;
assign p124 = c0;
assign p125 = c0;
assign p126 = c0;
assign p127 = c0;
assign p128 = c0;
assign p129 = c0;
assign p130 = c0;
assign p131 = c0;
assign p132 = c0;
assign p133 = c0;
assign p134 = c0;
assign p135 = c0;
assign p136 = c0;
assign p137 = c0;
assign p138 = c0;
assign p139 = c0;
assign p140 = c0;
assign p141 = c0;
assign p142 = c0;
assign p143 = c0;
assign p144 = c0;
assign p145 = c0;
assign p146 = c0;
assign p147 = c0;
assign p148 = c0;
assign p149 = c0;
assign p150 = c0;
assign p151 = c0;
assign p152 = c0;
assign p153 = c0;
assign p154 = c0;
assign p155 = c0;
assign p156 = c0;
assign p157 = c0;
assign p158 = c0;
assign p159 = c0;
assign p160 = c0;
assign p161 = c0;
assign p162 = c0;
assign p163 = c0;
assign p164 = c0;
assign p165 = c0;
assign p166 = c0;
assign p167 = c0;
assign p168 = c0;
assign p169 = c0;
assign p170 = c0;
assign p171 = c0;
assign p172 = c0;
assign p173 = c0;
assign p174 = c0;
assign p175 = c0;
assign p176 = c0;
assign p177 = c0;
assign p178 = c0;
assign p179 = c0;
assign p180 = c0;
assign p181 = c0;
assign p182 = c0;
assign p183 = c0;
assign p184 = c0;
assign p185 = c0;
assign p186 = c0;
assign p187 = c0;
assign p188 = c0;
assign p189 = c0;
assign p190 = c0;
assign p191 = c0;
assign p192 = c0;
assign p193 = c0;
assign p194 = c0;
assign p195 = c0;
assign p196 = c0;
assign p197 = c0;
assign p198 = c0;
assign p199 = c0;
assign p200 = c0;
assign p201 = c0;
assign p202 = c0;
assign p203 = c0;
assign p204 = c0;
assign p205 = c0;
assign p206 = c0;
assign p207 = c0;
assign p208 = c0;
assign p209 = c0;
assign p210 = c0;
assign p211 = c0;
assign p212 = c0;
assign p213 = c0;
assign p214 = c0;
assign p215 = c0;
assign p216 = c0;
assign p217 = c0;
assign p218 = c0;
assign p219 = c0;
assign p220 = c0;
assign p221 = c0;
assign p222 = c0;
assign p223 = c0;
assign p224 = c0;
assign p225 = c0;
assign p226 = c0;
assign p227 = c0;
assign p228 = c0;
assign p229 = c0;
assign p230 = c0;
assign p231 = c0;
assign p232 = c0;
assign p233 = c0;
assign p234 = c0;
assign p235 = c0;
assign p236 = c0;
assign p237 = c0;
assign p238 = c0;
assign p239 = c0;
assign p240 = c0;
assign p241 = c0;
assign p242 = c0;
assign p243 = c0;
assign p244 = c0;
assign p245 = c0;
assign p246 = c0;
assign p247 = c0;
assign p248 = c0;
assign p249 = c0;
assign p250 = c0;
assign p251 = c0;
assign p252 = c0;
assign p253 = c0;
assign p254 = c0;
assign p255 = c0;
assign p256 = c0;
assign p257 = c0;
assign p258 = c0;
assign p259 = c0;
assign p260 = c0;
assign p261 = c0;
assign p262 = c0;
assign p263 = c0;
assign p264 = c0;
assign p265 = c0;
assign p266 = c0;
assign p267 = c0;
assign p268 = c0;
assign p269 = c0;
assign p270 = c0;
assign p271 = c0;
assign p272 = c0;
assign p273 = c0;
assign p274 = c0;
assign p275 = c0;
assign p276 = c0;
assign p277 = c0;
assign p278 = c0;
assign p279 = c0;
assign p280 = c0;
assign p281 = c0;
assign p282 = c0;
assign p283 = c0;
assign p284 = c0;
assign p285 = c0;
assign p286 = c0;
assign p287 = c0;
assign p288 = c0;
assign p289 = c0;
assign p290 = c0;
assign p291 = c0;
assign p292 = c0;
assign p293 = c0;
assign p294 = c0;
assign p295 = c0;
assign p296 = c0;
assign p297 = c0;
assign p298 = c0;
assign p299 = c0;
assign p300 = c0;
assign p301 = c0;
assign p302 = c0;
assign p303 = c0;
assign p304 = c0;
assign p305 = c0;
assign p306 = c0;
assign p307 = c0;
assign p308 = c0;
assign p309 = c0;
assign p310 = c0;
assign p311 = c0;
assign p312 = c0;
assign p313 = c0;
assign p314 = c0;
assign p315 = c0;
assign p316 = c0;
assign p317 = c0;
assign p318 = c0;
assign p319 = c0;
assign p320 = c0;
assign p321 = c0;
assign p322 = c0;
assign p323 = c0;
assign p324 = c0;
assign p325 = c0;
assign p326 = c0;
assign p327 = c0;
assign p328 = c0;
assign p329 = c0;
assign p330 = c0;
assign p331 = c0;
assign p332 = c0;
assign p333 = c0;
assign p334 = c0;
assign p335 = c0;
assign p336 = c0;
assign p337 = c0;
assign p338 = c0;
assign p339 = c0;
assign p340 = c0;
assign p341 = c0;
assign p342 = c0;
assign p343 = c0;
assign p344 = c0;
assign p345 = c0;
assign p346 = c0;
assign p347 = c0;
assign p348 = c0;
assign p349 = c0;
assign p350 = c0;
assign p351 = c0;
assign p352 = c0;
assign p353 = c0;
assign p354 = c0;
assign p355 = c0;
assign p356 = c0;
assign p357 = c0;
assign p358 = c0;
assign p359 = c0;
assign p360 = c0;
assign p361 = c0;
assign p362 = c0;
assign p363 = c0;
assign p364 = c0;
assign p365 = c0;
assign p366 = c0;
assign p367 = c0;
assign p368 = c0;
assign p369 = c0;
assign p370 = c0;
assign p371 = c0;
assign p372 = c0;
assign p373 = c0;
assign p374 = c0;
assign p375 = c0;
assign p376 = c0;
assign p377 = c0;
assign p378 = c0;
assign p379 = c0;
assign p380 = c0;
assign p381 = c0;
assign p382 = c0;
assign p383 = c0;
assign p384 = c0;
assign p385 = c0;
assign p386 = c0;
assign p387 = c0;
assign p388 = c0;
assign p389 = c0;
assign p390 = c0;
assign p391 = c0;
assign p392 = c0;
assign p393 = c0;
assign p394 = c0;
assign p395 = c0;
assign p396 = c0;
assign p397 = c0;
assign p398 = c0;
assign p399 = c0;
assign p400 = c0;
assign p401 = c0;
assign p402 = c0;
assign p403 = c0;
assign p404 = c0;
assign p405 = c0;
assign p406 = c0;
assign p407 = c0;
assign p408 = c0;
assign p409 = c0;
assign p410 = c0;
assign p411 = c0;
assign p412 = c0;
assign p413 = c0;
assign p414 = c0;
assign p415 = c0;
assign p416 = c0;
assign p417 = c0;
assign p418 = c0;
assign p419 = c0;
assign p420 = c0;
assign p421 = c0;
assign p422 = c0;
assign p423 = c0;
assign p424 = c0;
assign p425 = c0;
assign p426 = c0;
assign p427 = c0;
assign p428 = c0;
assign p429 = c0;
assign p430 = c0;
assign p431 = c0;
assign p432 = c0;
assign p433 = c0;
assign p434 = c0;
assign p435 = c0;
assign p436 = c0;
assign p437 = c0;
assign p438 = c0;
assign p439 = c0;
assign p440 = c0;
assign p441 = c0;
assign p442 = c0;
assign p443 = c0;
assign p444 = c0;
assign p445 = c0;
assign p446 = c0;
assign p447 = c0;
assign p448 = c0;
assign p449 = c0;
assign p450 = c0;
assign p451 = c0;
assign p452 = c0;
assign p453 = c0;
assign p454 = c0;
assign p455 = c0;
assign p456 = c0;
assign p457 = c0;
assign p458 = c0;
assign p459 = c0;
assign p460 = c0;
assign p461 = c0;
assign p462 = c0;
assign p463 = c0;
assign p464 = c0;
assign p465 = c0;
assign p466 = c0;
assign p467 = c0;
assign p468 = c0;
assign p469 = c0;
assign p470 = c0;
assign p471 = c0;
assign p472 = c0;
assign p473 = c0;
assign p474 = c0;
assign p475 = c0;
assign p476 = c0;
assign p477 = c0;
assign p478 = c0;
assign p479 = c0;
assign p480 = c0;
assign p481 = c0;
assign p482 = c0;
assign p483 = c0;
assign p484 = c0;
assign p485 = c0;
assign p486 = c0;
assign p487 = c0;
assign p488 = c0;
assign p489 = c0;
assign p490 = c0;
assign p491 = c0;
assign p492 = c0;
assign p493 = c0;
assign p494 = c0;
assign p495 = c0;
assign p496 = c0;
assign p497 = c0;
assign p498 = c0;
assign p499 = c0;
assign p500 = c0;
assign p501 = c0;
assign p502 = c0;
assign p503 = c0;
assign p504 = c0;
assign p505 = c0;
assign p506 = c0;
assign p507 = c0;
assign p508 = c0;
assign p509 = c0;
assign p510 = c0;
assign p511 = c0;
assign p512 = c0;
assign p513 = c0;
assign p514 = c0;
assign p515 = c0;
assign p516 = c0;
assign p517 = c0;
assign p518 = c0;
assign p519 = c0;
assign p520 = c0;
assign p521 = c0;
assign p522 = c0;
assign p523 = c0;
assign p524 = c0;
assign p525 = c0;
assign p526 = c0;
assign p527 = c0;
assign p528 = c0;
assign p529 = c0;
assign p530 = c0;
assign p531 = c0;
assign p532 = c0;
assign p533 = c0;
assign p534 = c0;
assign p535 = c0;
assign p536 = c0;
assign p537 = c0;
assign p538 = c0;
assign p539 = c0;
assign p540 = c0;
assign p541 = c0;
assign p542 = c0;
assign p543 = c0;
assign p544 = c0;
assign p545 = c0;
assign p546 = c0;
assign p547 = c0;
assign p548 = c0;
assign p549 = c0;
assign p550 = c0;
assign p551 = c0;
assign p552 = c0;
assign p553 = c0;
assign p554 = c0;
assign p555 = c0;
assign p556 = c0;
assign p557 = c0;
assign p558 = c0;
assign p559 = c0;
assign p560 = c0;
assign p561 = c0;
assign p562 = c0;
assign p563 = c0;
assign p564 = c0;
assign p565 = c0;
assign p566 = c0;
assign p567 = c0;
assign p568 = c0;
assign p569 = c0;
assign p570 = c0;
assign p571 = c0;
assign p572 = c0;
assign p573 = c0;
assign p574 = c0;
assign p575 = c0;
assign p576 = c0;
assign p577 = c0;
assign p578 = c0;
assign p579 = c0;
assign p580 = c0;
assign p581 = c0;
assign p582 = c0;
assign p583 = c0;
assign p584 = c0;
assign p585 = c0;
assign p586 = c0;
assign p587 = c0;
assign p588 = c0;
assign p589 = c0;
assign p590 = c0;
assign p591 = c0;
assign p592 = c0;
assign p593 = c0;
assign p594 = c0;
assign p595 = c0;
assign p596 = c0;
assign p597 = c0;
assign p598 = c0;
assign p599 = c0;
assign p600 = c0;
assign p601 = c0;
assign p602 = c0;
assign p603 = c0;
assign p604 = c0;
assign p605 = c0;
assign p606 = c0;
assign p607 = c0;
assign p608 = c0;
assign p609 = c0;
assign p610 = c0;
assign p611 = c0;
assign p612 = c0;
assign p613 = c0;
assign p614 = c0;
assign p615 = c0;
assign p616 = c0;
assign p617 = c0;
assign p618 = c0;
assign p619 = c0;
assign p620 = c0;
assign p621 = c0;
assign p622 = c0;
assign p623 = c0;
assign p624 = c0;
assign p625 = c0;
assign p626 = c0;
assign p627 = c0;
assign p628 = c0;
assign p629 = c0;
assign p630 = c0;
assign p631 = c0;
assign p632 = c0;
assign p633 = c0;
assign p634 = c0;
assign p635 = c0;
assign p636 = c0;
assign p637 = c0;
assign p638 = c0;
assign p639 = c0;
assign p640 = c0;
assign p641 = c0;
assign p642 = c0;
assign p643 = c0;
assign p644 = c0;
assign p645 = c0;
assign p646 = c0;
assign p647 = c0;
assign p648 = c0;
assign p649 = c0;
assign p650 = c0;
assign p651 = c0;
assign p652 = c0;
assign p653 = c0;
assign p654 = c0;
assign p655 = c0;
assign p656 = c0;
assign p657 = c0;
assign p658 = c0;
assign p659 = c0;
assign p660 = c0;
assign p661 = c0;
assign p662 = c0;
assign p663 = c0;
assign p664 = c0;
assign p665 = c0;
assign p666 = c0;
assign p667 = c0;
assign p668 = c0;
assign p669 = c0;
assign p670 = c0;
assign p671 = c0;
assign p672 = c0;
assign p673 = c0;
assign p674 = c0;
assign p675 = c0;
assign p676 = c0;
assign p677 = c0;
assign p678 = c0;
assign p679 = c0;
assign p680 = c0;
assign p681 = c0;
assign p682 = c0;
assign p683 = c0;
assign p684 = c0;
assign p685 = c0;
assign p686 = c0;
assign p687 = c0;
assign p688 = c0;
assign p689 = c0;
assign p690 = c0;
assign p691 = c0;
assign p692 = c0;
assign p693 = c0;
assign p694 = c0;
assign p695 = c0;
assign p696 = c0;
assign p697 = c0;
assign p698 = c0;
assign p699 = c0;
assign p700 = c0;
assign p701 = c0;
assign p702 = c0;
assign p703 = c0;
assign p704 = c0;
assign p705 = c0;
assign p706 = c0;
assign p707 = c0;
assign p708 = c0;
assign p709 = c0;
assign p710 = c0;
assign p711 = c0;
assign p712 = c0;
assign p713 = c0;
assign p714 = c0;
assign p715 = c0;
assign p716 = c0;
assign p717 = c0;
assign p718 = c0;
assign p719 = c0;
assign p720 = c0;
assign p721 = c0;
assign p722 = c0;
assign p723 = c0;
assign p724 = c0;
assign p725 = c0;
assign p726 = c0;
assign p727 = c0;
assign p728 = c0;
assign p729 = c0;
assign p730 = c0;
assign p731 = c0;
assign p732 = c0;
assign p733 = c0;
assign p734 = c0;
assign p735 = c0;
assign p736 = c0;
assign p737 = c0;
assign p738 = c0;
assign p739 = c0;
assign p740 = c0;
assign p741 = c0;
assign p742 = c0;
assign p743 = c0;
assign p744 = c0;
assign p745 = c0;
assign p746 = c0;
assign p747 = c0;
assign p748 = c0;
assign p749 = c0;
assign p750 = c0;
assign p751 = c0;
assign p752 = c0;
assign p753 = c0;
assign p754 = c0;
assign p755 = c0;
assign p756 = c0;
assign p757 = c0;
assign p758 = c0;
assign p759 = c0;
assign p760 = c0;
assign p761 = c0;
assign p762 = c0;
assign p763 = c0;
assign p764 = c0;
assign p765 = c0;
assign p766 = c0;
assign p767 = c0;
assign p768 = c0;
assign p769 = c0;
assign p770 = c0;
assign p771 = c0;
assign p772 = c0;
assign p773 = c0;
assign p774 = c0;
assign p775 = c0;
assign p776 = c0;
assign p777 = c0;
assign p778 = c0;
assign p779 = c0;
assign p780 = c0;
assign p781 = c0;
assign p782 = c0;
assign p783 = c0;
assign p784 = c0;
assign p785 = c0;
assign p786 = c0;
assign p787 = c0;
assign p788 = c0;
assign p789 = c0;
assign p790 = c0;
assign p791 = c0;
assign p792 = c0;
assign p793 = c0;
assign p794 = c0;
assign p795 = c0;
assign p796 = c0;
assign p797 = c0;
assign p798 = c0;
assign p799 = c0;
assign p800 = c0;
assign p801 = c0;
assign p802 = c0;
assign p803 = c0;
assign p804 = c0;
assign p805 = c0;
assign p806 = c0;
assign p807 = c0;
assign p808 = c0;
assign p809 = c0;
assign p810 = c0;
assign p811 = c0;
assign p812 = c0;
assign p813 = c0;
assign p814 = c0;
assign p815 = c0;
assign p816 = c0;
assign p817 = c0;
assign p818 = c0;
assign p819 = c0;
assign p820 = c0;
assign p821 = c0;
assign p822 = c0;
assign p823 = c0;
assign p824 = c0;
assign p825 = c0;
assign p826 = c0;
assign p827 = c0;
assign p828 = c0;
assign p829 = c0;
assign p830 = c0;
assign p831 = c0;
assign p832 = c0;
assign p833 = c0;
assign p834 = c0;
assign p835 = c0;
assign p836 = c0;
assign p837 = c0;
assign p838 = c0;
assign p839 = c0;
assign p840 = c0;
assign p841 = c0;
assign p842 = c0;
assign p843 = c0;
assign p844 = c0;
assign p845 = c0;
assign p846 = c0;
assign p847 = c0;
assign p848 = c0;
assign p849 = c0;
assign p850 = c0;
assign p851 = c0;
assign p852 = c0;
assign p853 = c0;
assign p854 = c0;
assign p855 = c0;
assign p856 = c0;
assign p857 = c0;
assign p858 = c0;
assign p859 = c0;
assign p860 = c0;
assign p861 = c0;
assign p862 = c0;
assign p863 = c0;
assign p864 = c0;
assign p865 = c0;
assign p866 = c0;
assign p867 = c0;
assign p868 = c0;
assign p869 = c0;
assign p870 = c0;
assign p871 = c0;
assign p872 = c0;
assign p873 = c0;
assign p874 = c0;
assign p875 = c0;
assign p876 = c0;
assign p877 = c0;
assign p878 = c0;
assign p879 = c0;
assign p880 = c0;
assign p881 = c0;
assign p882 = c0;
assign p883 = c0;
assign p884 = c0;
assign p885 = c0;
assign p886 = c0;
assign p887 = c0;
assign p888 = c0;
assign p889 = c0;
assign p890 = c0;
assign p891 = c0;
assign p892 = c0;
assign p893 = c0;
assign p894 = c0;
assign p895 = c0;
assign p896 = c0;
assign p897 = c0;
assign p898 = c0;
assign p899 = c0;
assign p900 = c0;
assign p901 = c0;
assign p902 = c0;
assign p903 = c0;
assign p904 = c0;
assign p905 = c0;
assign p906 = c0;
assign p907 = c0;
assign p908 = c0;
assign p909 = c0;
assign p910 = c0;
assign p911 = c0;
assign p912 = c0;
assign p913 = c0;
assign p914 = c0;
assign p915 = c0;
assign p916 = c0;
assign p917 = c0;
assign p918 = c0;
assign p919 = c0;
assign p920 = c0;
assign p921 = c0;
assign p922 = c0;
assign p923 = c0;
assign p924 = c0;
assign p925 = c0;
assign p926 = c0;
assign p927 = l994;
assign p928 = c0;
assign p929 = c0;
assign p930 = a1024;
assign p931 = c0;
assign p932 = c0;
assign p933 = a1032;
assign p934 = a1040;
assign p935 = a1046;
assign p936 = a1052;
assign p937 = a1056;
assign p938 = a1060;
assign p939 = a1064;
assign p940 = a1068;
assign p941 = a1076;
assign p942 = a1080;
assign p943 = a1082;
assign p944 = a1096;
assign p945 = a1100;
assign p946 = a1104;
assign p947 = a1106;
assign p948 = a1236;
assign p949 = a1248;
assign p950 = a1252;
assign p951 = ~a1258;
assign p952 = ~a1274;
assign p953 = a1296;
assign p954 = a1320;
assign p955 = c0;
assign p956 = c0;
assign p957 = c0;
assign p958 = c0;
assign p959 = c0;
assign p960 = c0;
assign p961 = c0;
assign p962 = c0;
assign p963 = c0;
assign p964 = c0;
assign p965 = c0;
assign p966 = c0;
assign p967 = c0;
assign p968 = c0;
assign p969 = c0;
assign p970 = c0;
assign p971 = c0;
assign p972 = c0;
assign p973 = c0;
assign p974 = c0;
assign p975 = c0;
assign p976 = c0;
assign p977 = c0;
assign p978 = c0;
assign p979 = c0;
assign p980 = c0;
assign p981 = c0;
assign p982 = c0;
assign p983 = c0;
assign p984 = c0;
assign p985 = c0;
assign p986 = c0;
assign p987 = c0;
assign p988 = c0;
assign p989 = c0;
assign p990 = c0;
assign p991 = c0;
assign p992 = c0;
assign p993 = c0;
assign p994 = c0;
assign p995 = c0;
assign p996 = c0;
assign p997 = c0;
assign p998 = c0;
assign p999 = c0;
assign p1000 = c0;
assign p1001 = c0;
assign p1002 = c0;
assign p1003 = c0;
assign p1004 = c0;
assign p1005 = c0;
assign p1006 = c0;
assign p1007 = c0;
assign p1008 = c0;
assign p1009 = c0;
assign p1010 = c0;
assign p1011 = c0;
assign p1012 = c0;
assign p1013 = c0;
assign p1014 = c0;
assign p1015 = c0;
assign p1016 = a1322;
assign p1017 = a1360;
assign p1018 = a1368;
assign p1019 = a1378;
assign p1020 = a1352;
assign p1021 = a1388;
assign p1022 = a1404;
assign p1023 = ~a1426;
assign p1024 = c0;
assign p1025 = a1476;
assign p1026 = ~a1482;
assign p1027 = a1486;
assign p1028 = ~a1494;
assign p1029 = a1506;
assign p1030 = a1588;
assign p1031 = a1660;
assign p1032 = a1664;
assign p1033 = a1668;
assign p1034 = c0;
assign p1035 = a1702;
assign p1036 = a2308;
assign p1037 = c0;
assign p1038 = ~a2382;
assign p1039 = c0;
assign p1040 = c0;
assign p1041 = c0;
assign p1042 = ~a2456;
assign p1043 = a2458;
assign p1044 = ~a2460;
assign p1045 = c0;
assign p1046 = ~a2530;
assign p1047 = a2532;
assign p1048 = a2534;
assign p1049 = ~a2536;
assign p1050 = c0;
assign p1051 = c0;
assign p1052 = c0;
assign p1053 = c0;
assign p1054 = c0;
assign p1055 = c0;
assign p1056 = c0;
assign p1057 = c0;
assign p1058 = c0;
assign p1059 = c0;
assign p1060 = c0;
assign p1061 = c0;
assign p1062 = c0;
assign p1063 = c0;
assign p1064 = c0;
assign p1065 = c0;
assign p1066 = c0;
assign p1067 = c0;
assign p1068 = c0;
assign p1069 = c0;
assign p1070 = c0;
assign p1071 = c0;
assign p1072 = c0;
assign p1073 = c0;
assign p1074 = c0;
assign p1075 = c0;
assign p1076 = c0;
assign p1077 = c0;
assign p1078 = c0;
assign p1079 = a2544;
assign p1080 = c0;
assign p1081 = c0;
assign p1082 = c0;
assign p1083 = c0;
assign p1084 = c0;
assign p1085 = c0;
assign p1086 = c0;
assign p1087 = c0;
assign p1088 = c0;
assign p1089 = c0;
assign p1090 = c0;
assign p1091 = c0;
assign p1092 = c0;
assign p1093 = c0;
assign p1094 = c0;
assign p1095 = c0;
assign p1096 = c0;
assign p1097 = c0;
assign p1098 = c0;
assign p1099 = c0;
assign p1100 = c0;
assign p1101 = c0;
assign p1102 = c0;
assign p1103 = c0;
assign p1104 = c0;
assign p1105 = c0;
assign p1106 = c0;
assign p1107 = c0;
assign p1108 = c0;
assign p1109 = c0;
assign p1110 = c0;
assign p1111 = c0;
assign p1112 = c0;
assign p1113 = c0;
assign p1114 = c0;
assign p1115 = c0;
assign p1116 = c0;
assign p1117 = c0;
assign p1118 = c0;
assign p1119 = c0;
assign p1120 = c0;
assign p1121 = c0;
assign p1122 = c0;
assign p1123 = c0;
assign p1124 = c0;
assign p1125 = c0;
assign p1126 = c0;
assign p1127 = c0;
assign p1128 = c0;
assign p1129 = c0;
assign p1130 = c0;
assign p1131 = c0;
assign p1132 = c0;
assign p1133 = c0;
assign p1134 = c0;
assign p1135 = c0;
assign p1136 = c0;
assign p1137 = a2590;
assign p1138 = a2636;
assign p1139 = c0;
assign p1140 = c0;
assign p1141 = c0;
assign p1142 = a2544;
assign p1143 = c0;
assign p1144 = a2650;
assign p1145 = c0;
assign p1146 = c0;
assign p1147 = c0;
assign p1148 = a2676;
assign p1149 = a2690;

assert property (~p0);
assert property (~p1);
assert property (~p2);
assert property (~p3);
assert property (~p4);
assert property (~p5);
assert property (~p6);
assert property (~p7);
assert property (~p8);
assert property (~p9);
assert property (~p10);
assert property (~p11);
assert property (~p12);
assert property (~p13);
assert property (~p14);
assert property (~p15);
assert property (~p16);
assert property (~p17);
assert property (~p18);
assert property (~p19);
assert property (~p20);
assert property (~p21);
assert property (~p22);
assert property (~p23);
assert property (~p24);
assert property (~p25);
assert property (~p26);
assert property (~p27);
assert property (~p28);
assert property (~p29);
assert property (~p30);
assert property (~p31);
assert property (~p32);
assert property (~p33);
assert property (~p34);
assert property (~p35);
assert property (~p36);
assert property (~p37);
assert property (~p38);
assert property (~p39);
assert property (~p40);
assert property (~p41);
assert property (~p42);
assert property (~p43);
assert property (~p44);
assert property (~p45);
assert property (~p46);
assert property (~p47);
assert property (~p48);
assert property (~p49);
assert property (~p50);
assert property (~p51);
assert property (~p52);
assert property (~p53);
assert property (~p54);
assert property (~p55);
assert property (~p56);
assert property (~p57);
assert property (~p58);
assert property (~p59);
assert property (~p60);
assert property (~p61);
assert property (~p62);
assert property (~p63);
assert property (~p64);
assert property (~p65);
assert property (~p66);
assert property (~p67);
assert property (~p68);
assert property (~p69);
assert property (~p70);
assert property (~p71);
assert property (~p72);
assert property (~p73);
assert property (~p74);
assert property (~p75);
assert property (~p76);
assert property (~p77);
assert property (~p78);
assert property (~p79);
assert property (~p80);
assert property (~p81);
assert property (~p82);
assert property (~p83);
assert property (~p84);
assert property (~p85);
assert property (~p86);
assert property (~p87);
assert property (~p88);
assert property (~p89);
assert property (~p90);
assert property (~p91);
assert property (~p92);
assert property (~p93);
assert property (~p94);
assert property (~p95);
assert property (~p96);
assert property (~p97);
assert property (~p98);
assert property (~p99);
assert property (~p100);
assert property (~p101);
assert property (~p102);
assert property (~p103);
assert property (~p104);
assert property (~p105);
assert property (~p106);
assert property (~p107);
assert property (~p108);
assert property (~p109);
assert property (~p110);
assert property (~p111);
assert property (~p112);
assert property (~p113);
assert property (~p114);
assert property (~p115);
assert property (~p116);
assert property (~p117);
assert property (~p118);
assert property (~p119);
assert property (~p120);
assert property (~p121);
assert property (~p122);
assert property (~p123);
assert property (~p124);
assert property (~p125);
assert property (~p126);
assert property (~p127);
assert property (~p128);
assert property (~p129);
assert property (~p130);
assert property (~p131);
assert property (~p132);
assert property (~p133);
assert property (~p134);
assert property (~p135);
assert property (~p136);
assert property (~p137);
assert property (~p138);
assert property (~p139);
assert property (~p140);
assert property (~p141);
assert property (~p142);
assert property (~p143);
assert property (~p144);
assert property (~p145);
assert property (~p146);
assert property (~p147);
assert property (~p148);
assert property (~p149);
assert property (~p150);
assert property (~p151);
assert property (~p152);
assert property (~p153);
assert property (~p154);
assert property (~p155);
assert property (~p156);
assert property (~p157);
assert property (~p158);
assert property (~p159);
assert property (~p160);
assert property (~p161);
assert property (~p162);
assert property (~p163);
assert property (~p164);
assert property (~p165);
assert property (~p166);
assert property (~p167);
assert property (~p168);
assert property (~p169);
assert property (~p170);
assert property (~p171);
assert property (~p172);
assert property (~p173);
assert property (~p174);
assert property (~p175);
assert property (~p176);
assert property (~p177);
assert property (~p178);
assert property (~p179);
assert property (~p180);
assert property (~p181);
assert property (~p182);
assert property (~p183);
assert property (~p184);
assert property (~p185);
assert property (~p186);
assert property (~p187);
assert property (~p188);
assert property (~p189);
assert property (~p190);
assert property (~p191);
assert property (~p192);
assert property (~p193);
assert property (~p194);
assert property (~p195);
assert property (~p196);
assert property (~p197);
assert property (~p198);
assert property (~p199);
assert property (~p200);
assert property (~p201);
assert property (~p202);
assert property (~p203);
assert property (~p204);
assert property (~p205);
assert property (~p206);
assert property (~p207);
assert property (~p208);
assert property (~p209);
assert property (~p210);
assert property (~p211);
assert property (~p212);
assert property (~p213);
assert property (~p214);
assert property (~p215);
assert property (~p216);
assert property (~p217);
assert property (~p218);
assert property (~p219);
assert property (~p220);
assert property (~p221);
assert property (~p222);
assert property (~p223);
assert property (~p224);
assert property (~p225);
assert property (~p226);
assert property (~p227);
assert property (~p228);
assert property (~p229);
assert property (~p230);
assert property (~p231);
assert property (~p232);
assert property (~p233);
assert property (~p234);
assert property (~p235);
assert property (~p236);
assert property (~p237);
assert property (~p238);
assert property (~p239);
assert property (~p240);
assert property (~p241);
assert property (~p242);
assert property (~p243);
assert property (~p244);
assert property (~p245);
assert property (~p246);
assert property (~p247);
assert property (~p248);
assert property (~p249);
assert property (~p250);
assert property (~p251);
assert property (~p252);
assert property (~p253);
assert property (~p254);
assert property (~p255);
assert property (~p256);
assert property (~p257);
assert property (~p258);
assert property (~p259);
assert property (~p260);
assert property (~p261);
assert property (~p262);
assert property (~p263);
assert property (~p264);
assert property (~p265);
assert property (~p266);
assert property (~p267);
assert property (~p268);
assert property (~p269);
assert property (~p270);
assert property (~p271);
assert property (~p272);
assert property (~p273);
assert property (~p274);
assert property (~p275);
assert property (~p276);
assert property (~p277);
assert property (~p278);
assert property (~p279);
assert property (~p280);
assert property (~p281);
assert property (~p282);
assert property (~p283);
assert property (~p284);
assert property (~p285);
assert property (~p286);
assert property (~p287);
assert property (~p288);
assert property (~p289);
assert property (~p290);
assert property (~p291);
assert property (~p292);
assert property (~p293);
assert property (~p294);
assert property (~p295);
assert property (~p296);
assert property (~p297);
assert property (~p298);
assert property (~p299);
assert property (~p300);
assert property (~p301);
assert property (~p302);
assert property (~p303);
assert property (~p304);
assert property (~p305);
assert property (~p306);
assert property (~p307);
assert property (~p308);
assert property (~p309);
assert property (~p310);
assert property (~p311);
assert property (~p312);
assert property (~p313);
assert property (~p314);
assert property (~p315);
assert property (~p316);
assert property (~p317);
assert property (~p318);
assert property (~p319);
assert property (~p320);
assert property (~p321);
assert property (~p322);
assert property (~p323);
assert property (~p324);
assert property (~p325);
assert property (~p326);
assert property (~p327);
assert property (~p328);
assert property (~p329);
assert property (~p330);
assert property (~p331);
assert property (~p332);
assert property (~p333);
assert property (~p334);
assert property (~p335);
assert property (~p336);
assert property (~p337);
assert property (~p338);
assert property (~p339);
assert property (~p340);
assert property (~p341);
assert property (~p342);
assert property (~p343);
assert property (~p344);
assert property (~p345);
assert property (~p346);
assert property (~p347);
assert property (~p348);
assert property (~p349);
assert property (~p350);
assert property (~p351);
assert property (~p352);
assert property (~p353);
assert property (~p354);
assert property (~p355);
assert property (~p356);
assert property (~p357);
assert property (~p358);
assert property (~p359);
assert property (~p360);
assert property (~p361);
assert property (~p362);
assert property (~p363);
assert property (~p364);
assert property (~p365);
assert property (~p366);
assert property (~p367);
assert property (~p368);
assert property (~p369);
assert property (~p370);
assert property (~p371);
assert property (~p372);
assert property (~p373);
assert property (~p374);
assert property (~p375);
assert property (~p376);
assert property (~p377);
assert property (~p378);
assert property (~p379);
assert property (~p380);
assert property (~p381);
assert property (~p382);
assert property (~p383);
assert property (~p384);
assert property (~p385);
assert property (~p386);
assert property (~p387);
assert property (~p388);
assert property (~p389);
assert property (~p390);
assert property (~p391);
assert property (~p392);
assert property (~p393);
assert property (~p394);
assert property (~p395);
assert property (~p396);
assert property (~p397);
assert property (~p398);
assert property (~p399);
assert property (~p400);
assert property (~p401);
assert property (~p402);
assert property (~p403);
assert property (~p404);
assert property (~p405);
assert property (~p406);
assert property (~p407);
assert property (~p408);
assert property (~p409);
assert property (~p410);
assert property (~p411);
assert property (~p412);
assert property (~p413);
assert property (~p414);
assert property (~p415);
assert property (~p416);
assert property (~p417);
assert property (~p418);
assert property (~p419);
assert property (~p420);
assert property (~p421);
assert property (~p422);
assert property (~p423);
assert property (~p424);
assert property (~p425);
assert property (~p426);
assert property (~p427);
assert property (~p428);
assert property (~p429);
assert property (~p430);
assert property (~p431);
assert property (~p432);
assert property (~p433);
assert property (~p434);
assert property (~p435);
assert property (~p436);
assert property (~p437);
assert property (~p438);
assert property (~p439);
assert property (~p440);
assert property (~p441);
assert property (~p442);
assert property (~p443);
assert property (~p444);
assert property (~p445);
assert property (~p446);
assert property (~p447);
assert property (~p448);
assert property (~p449);
assert property (~p450);
assert property (~p451);
assert property (~p452);
assert property (~p453);
assert property (~p454);
assert property (~p455);
assert property (~p456);
assert property (~p457);
assert property (~p458);
assert property (~p459);
assert property (~p460);
assert property (~p461);
assert property (~p462);
assert property (~p463);
assert property (~p464);
assert property (~p465);
assert property (~p466);
assert property (~p467);
assert property (~p468);
assert property (~p469);
assert property (~p470);
assert property (~p471);
assert property (~p472);
assert property (~p473);
assert property (~p474);
assert property (~p475);
assert property (~p476);
assert property (~p477);
assert property (~p478);
assert property (~p479);
assert property (~p480);
assert property (~p481);
assert property (~p482);
assert property (~p483);
assert property (~p484);
assert property (~p485);
assert property (~p486);
assert property (~p487);
assert property (~p488);
assert property (~p489);
assert property (~p490);
assert property (~p491);
assert property (~p492);
assert property (~p493);
assert property (~p494);
assert property (~p495);
assert property (~p496);
assert property (~p497);
assert property (~p498);
assert property (~p499);
assert property (~p500);
assert property (~p501);
assert property (~p502);
assert property (~p503);
assert property (~p504);
assert property (~p505);
assert property (~p506);
assert property (~p507);
assert property (~p508);
assert property (~p509);
assert property (~p510);
assert property (~p511);
assert property (~p512);
assert property (~p513);
assert property (~p514);
assert property (~p515);
assert property (~p516);
assert property (~p517);
assert property (~p518);
assert property (~p519);
assert property (~p520);
assert property (~p521);
assert property (~p522);
assert property (~p523);
assert property (~p524);
assert property (~p525);
assert property (~p526);
assert property (~p527);
assert property (~p528);
assert property (~p529);
assert property (~p530);
assert property (~p531);
assert property (~p532);
assert property (~p533);
assert property (~p534);
assert property (~p535);
assert property (~p536);
assert property (~p537);
assert property (~p538);
assert property (~p539);
assert property (~p540);
assert property (~p541);
assert property (~p542);
assert property (~p543);
assert property (~p544);
assert property (~p545);
assert property (~p546);
assert property (~p547);
assert property (~p548);
assert property (~p549);
assert property (~p550);
assert property (~p551);
assert property (~p552);
assert property (~p553);
assert property (~p554);
assert property (~p555);
assert property (~p556);
assert property (~p557);
assert property (~p558);
assert property (~p559);
assert property (~p560);
assert property (~p561);
assert property (~p562);
assert property (~p563);
assert property (~p564);
assert property (~p565);
assert property (~p566);
assert property (~p567);
assert property (~p568);
assert property (~p569);
assert property (~p570);
assert property (~p571);
assert property (~p572);
assert property (~p573);
assert property (~p574);
assert property (~p575);
assert property (~p576);
assert property (~p577);
assert property (~p578);
assert property (~p579);
assert property (~p580);
assert property (~p581);
assert property (~p582);
assert property (~p583);
assert property (~p584);
assert property (~p585);
assert property (~p586);
assert property (~p587);
assert property (~p588);
assert property (~p589);
assert property (~p590);
assert property (~p591);
assert property (~p592);
assert property (~p593);
assert property (~p594);
assert property (~p595);
assert property (~p596);
assert property (~p597);
assert property (~p598);
assert property (~p599);
assert property (~p600);
assert property (~p601);
assert property (~p602);
assert property (~p603);
assert property (~p604);
assert property (~p605);
assert property (~p606);
assert property (~p607);
assert property (~p608);
assert property (~p609);
assert property (~p610);
assert property (~p611);
assert property (~p612);
assert property (~p613);
assert property (~p614);
assert property (~p615);
assert property (~p616);
assert property (~p617);
assert property (~p618);
assert property (~p619);
assert property (~p620);
assert property (~p621);
assert property (~p622);
assert property (~p623);
assert property (~p624);
assert property (~p625);
assert property (~p626);
assert property (~p627);
assert property (~p628);
assert property (~p629);
assert property (~p630);
assert property (~p631);
assert property (~p632);
assert property (~p633);
assert property (~p634);
assert property (~p635);
assert property (~p636);
assert property (~p637);
assert property (~p638);
assert property (~p639);
assert property (~p640);
assert property (~p641);
assert property (~p642);
assert property (~p643);
assert property (~p644);
assert property (~p645);
assert property (~p646);
assert property (~p647);
assert property (~p648);
assert property (~p649);
assert property (~p650);
assert property (~p651);
assert property (~p652);
assert property (~p653);
assert property (~p654);
assert property (~p655);
assert property (~p656);
assert property (~p657);
assert property (~p658);
assert property (~p659);
assert property (~p660);
assert property (~p661);
assert property (~p662);
assert property (~p663);
assert property (~p664);
assert property (~p665);
assert property (~p666);
assert property (~p667);
assert property (~p668);
assert property (~p669);
assert property (~p670);
assert property (~p671);
assert property (~p672);
assert property (~p673);
assert property (~p674);
assert property (~p675);
assert property (~p676);
assert property (~p677);
assert property (~p678);
assert property (~p679);
assert property (~p680);
assert property (~p681);
assert property (~p682);
assert property (~p683);
assert property (~p684);
assert property (~p685);
assert property (~p686);
assert property (~p687);
assert property (~p688);
assert property (~p689);
assert property (~p690);
assert property (~p691);
assert property (~p692);
assert property (~p693);
assert property (~p694);
assert property (~p695);
assert property (~p696);
assert property (~p697);
assert property (~p698);
assert property (~p699);
assert property (~p700);
assert property (~p701);
assert property (~p702);
assert property (~p703);
assert property (~p704);
assert property (~p705);
assert property (~p706);
assert property (~p707);
assert property (~p708);
assert property (~p709);
assert property (~p710);
assert property (~p711);
assert property (~p712);
assert property (~p713);
assert property (~p714);
assert property (~p715);
assert property (~p716);
assert property (~p717);
assert property (~p718);
assert property (~p719);
assert property (~p720);
assert property (~p721);
assert property (~p722);
assert property (~p723);
assert property (~p724);
assert property (~p725);
assert property (~p726);
assert property (~p727);
assert property (~p728);
assert property (~p729);
assert property (~p730);
assert property (~p731);
assert property (~p732);
assert property (~p733);
assert property (~p734);
assert property (~p735);
assert property (~p736);
assert property (~p737);
assert property (~p738);
assert property (~p739);
assert property (~p740);
assert property (~p741);
assert property (~p742);
assert property (~p743);
assert property (~p744);
assert property (~p745);
assert property (~p746);
assert property (~p747);
assert property (~p748);
assert property (~p749);
assert property (~p750);
assert property (~p751);
assert property (~p752);
assert property (~p753);
assert property (~p754);
assert property (~p755);
assert property (~p756);
assert property (~p757);
assert property (~p758);
assert property (~p759);
assert property (~p760);
assert property (~p761);
assert property (~p762);
assert property (~p763);
assert property (~p764);
assert property (~p765);
assert property (~p766);
assert property (~p767);
assert property (~p768);
assert property (~p769);
assert property (~p770);
assert property (~p771);
assert property (~p772);
assert property (~p773);
assert property (~p774);
assert property (~p775);
assert property (~p776);
assert property (~p777);
assert property (~p778);
assert property (~p779);
assert property (~p780);
assert property (~p781);
assert property (~p782);
assert property (~p783);
assert property (~p784);
assert property (~p785);
assert property (~p786);
assert property (~p787);
assert property (~p788);
assert property (~p789);
assert property (~p790);
assert property (~p791);
assert property (~p792);
assert property (~p793);
assert property (~p794);
assert property (~p795);
assert property (~p796);
assert property (~p797);
assert property (~p798);
assert property (~p799);
assert property (~p800);
assert property (~p801);
assert property (~p802);
assert property (~p803);
assert property (~p804);
assert property (~p805);
assert property (~p806);
assert property (~p807);
assert property (~p808);
assert property (~p809);
assert property (~p810);
assert property (~p811);
assert property (~p812);
assert property (~p813);
assert property (~p814);
assert property (~p815);
assert property (~p816);
assert property (~p817);
assert property (~p818);
assert property (~p819);
assert property (~p820);
assert property (~p821);
assert property (~p822);
assert property (~p823);
assert property (~p824);
assert property (~p825);
assert property (~p826);
assert property (~p827);
assert property (~p828);
assert property (~p829);
assert property (~p830);
assert property (~p831);
assert property (~p832);
assert property (~p833);
assert property (~p834);
assert property (~p835);
assert property (~p836);
assert property (~p837);
assert property (~p838);
assert property (~p839);
assert property (~p840);
assert property (~p841);
assert property (~p842);
assert property (~p843);
assert property (~p844);
assert property (~p845);
assert property (~p846);
assert property (~p847);
assert property (~p848);
assert property (~p849);
assert property (~p850);
assert property (~p851);
assert property (~p852);
assert property (~p853);
assert property (~p854);
assert property (~p855);
assert property (~p856);
assert property (~p857);
assert property (~p858);
assert property (~p859);
assert property (~p860);
assert property (~p861);
assert property (~p862);
assert property (~p863);
assert property (~p864);
assert property (~p865);
assert property (~p866);
assert property (~p867);
assert property (~p868);
assert property (~p869);
assert property (~p870);
assert property (~p871);
assert property (~p872);
assert property (~p873);
assert property (~p874);
assert property (~p875);
assert property (~p876);
assert property (~p877);
assert property (~p878);
assert property (~p879);
assert property (~p880);
assert property (~p881);
assert property (~p882);
assert property (~p883);
assert property (~p884);
assert property (~p885);
assert property (~p886);
assert property (~p887);
assert property (~p888);
assert property (~p889);
assert property (~p890);
assert property (~p891);
assert property (~p892);
assert property (~p893);
assert property (~p894);
assert property (~p895);
assert property (~p896);
assert property (~p897);
assert property (~p898);
assert property (~p899);
assert property (~p900);
assert property (~p901);
assert property (~p902);
assert property (~p903);
assert property (~p904);
assert property (~p905);
assert property (~p906);
assert property (~p907);
assert property (~p908);
assert property (~p909);
assert property (~p910);
assert property (~p911);
assert property (~p912);
assert property (~p913);
assert property (~p914);
assert property (~p915);
assert property (~p916);
assert property (~p917);
assert property (~p918);
assert property (~p919);
assert property (~p920);
assert property (~p921);
assert property (~p922);
assert property (~p923);
assert property (~p924);
assert property (~p925);
assert property (~p926);
assert property (~p927);
assert property (~p928);
assert property (~p929);
assert property (~p930);
assert property (~p931);
assert property (~p932);
assert property (~p933);
assert property (~p934);
assert property (~p935);
assert property (~p936);
assert property (~p937);
assert property (~p938);
assert property (~p939);
assert property (~p940);
assert property (~p941);
assert property (~p942);
assert property (~p943);
assert property (~p944);
assert property (~p945);
assert property (~p946);
assert property (~p947);
assert property (~p948);
assert property (~p949);
assert property (~p950);
assert property (~p951);
assert property (~p952);
assert property (~p953);
assert property (~p954);
assert property (~p955);
assert property (~p956);
assert property (~p957);
assert property (~p958);
assert property (~p959);
assert property (~p960);
assert property (~p961);
assert property (~p962);
assert property (~p963);
assert property (~p964);
assert property (~p965);
assert property (~p966);
assert property (~p967);
assert property (~p968);
assert property (~p969);
assert property (~p970);
assert property (~p971);
assert property (~p972);
assert property (~p973);
assert property (~p974);
assert property (~p975);
assert property (~p976);
assert property (~p977);
assert property (~p978);
assert property (~p979);
assert property (~p980);
assert property (~p981);
assert property (~p982);
assert property (~p983);
assert property (~p984);
assert property (~p985);
assert property (~p986);
assert property (~p987);
assert property (~p988);
assert property (~p989);
assert property (~p990);
assert property (~p991);
assert property (~p992);
assert property (~p993);
assert property (~p994);
assert property (~p995);
assert property (~p996);
assert property (~p997);
assert property (~p998);
assert property (~p999);
assert property (~p1000);
assert property (~p1001);
assert property (~p1002);
assert property (~p1003);
assert property (~p1004);
assert property (~p1005);
assert property (~p1006);
assert property (~p1007);
assert property (~p1008);
assert property (~p1009);
assert property (~p1010);
assert property (~p1011);
assert property (~p1012);
assert property (~p1013);
assert property (~p1014);
assert property (~p1015);
assert property (~p1016);
assert property (~p1017);
assert property (~p1018);
assert property (~p1019);
assert property (~p1020);
assert property (~p1021);
assert property (~p1022);
assert property (~p1023);
assert property (~p1024);
assert property (~p1025);
assert property (~p1026);
assert property (~p1027);
assert property (~p1028);
assert property (~p1029);
assert property (~p1030);
assert property (~p1031);
assert property (~p1032);
assert property (~p1033);
assert property (~p1034);
assert property (~p1035);
assert property (~p1036);
assert property (~p1037);
assert property (~p1038);
assert property (~p1039);
assert property (~p1040);
assert property (~p1041);
assert property (~p1042);
assert property (~p1043);
assert property (~p1044);
assert property (~p1045);
assert property (~p1046);
assert property (~p1047);
assert property (~p1048);
assert property (~p1049);
assert property (~p1050);
assert property (~p1051);
assert property (~p1052);
assert property (~p1053);
assert property (~p1054);
assert property (~p1055);
assert property (~p1056);
assert property (~p1057);
assert property (~p1058);
assert property (~p1059);
assert property (~p1060);
assert property (~p1061);
assert property (~p1062);
assert property (~p1063);
assert property (~p1064);
assert property (~p1065);
assert property (~p1066);
assert property (~p1067);
assert property (~p1068);
assert property (~p1069);
assert property (~p1070);
assert property (~p1071);
assert property (~p1072);
assert property (~p1073);
assert property (~p1074);
assert property (~p1075);
assert property (~p1076);
assert property (~p1077);
assert property (~p1078);
assert property (~p1079);
assert property (~p1080);
assert property (~p1081);
assert property (~p1082);
assert property (~p1083);
assert property (~p1084);
assert property (~p1085);
assert property (~p1086);
assert property (~p1087);
assert property (~p1088);
assert property (~p1089);
assert property (~p1090);
assert property (~p1091);
assert property (~p1092);
assert property (~p1093);
assert property (~p1094);
assert property (~p1095);
assert property (~p1096);
assert property (~p1097);
assert property (~p1098);
assert property (~p1099);
assert property (~p1100);
assert property (~p1101);
assert property (~p1102);
assert property (~p1103);
assert property (~p1104);
assert property (~p1105);
assert property (~p1106);
assert property (~p1107);
assert property (~p1108);
assert property (~p1109);
assert property (~p1110);
assert property (~p1111);
assert property (~p1112);
assert property (~p1113);
assert property (~p1114);
assert property (~p1115);
assert property (~p1116);
assert property (~p1117);
assert property (~p1118);
assert property (~p1119);
assert property (~p1120);
assert property (~p1121);
assert property (~p1122);
assert property (~p1123);
assert property (~p1124);
assert property (~p1125);
assert property (~p1126);
assert property (~p1127);
assert property (~p1128);
assert property (~p1129);
assert property (~p1130);
assert property (~p1131);
assert property (~p1132);
assert property (~p1133);
assert property (~p1134);
assert property (~p1135);
assert property (~p1136);
assert property (~p1137);
assert property (~p1138);
assert property (~p1139);
assert property (~p1140);
assert property (~p1141);
assert property (~p1142);
assert property (~p1143);
assert property (~p1144);
assert property (~p1145);
assert property (~p1146);
assert property (~p1147);
assert property (~p1148);
assert property (~p1149);

endmodule
