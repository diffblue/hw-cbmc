module main;

  // === takes any type except real/shortreal
  wire x = 1.1 === 1.2;

endmodule
