// as 'description'
typedef bit my_type1;

module main();

  // as 'module_item'
  typedef bit my_type2;

  function some_function;
    // as 'block_item'
    typedef bit my_type3;
    begin
    end
  endfunction

endmodule
