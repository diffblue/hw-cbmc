checker myChecker;
endchecker

module main;
endmodule
