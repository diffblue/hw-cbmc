module pdtvispeterson (i2,i4,p0);

input i2,i4;

output p0;

wire na162,na228,na776,na800,na822,na1334,na1358,na1380,na1424,a26,a28,a30,a32,a34,a36,
a38,a40,a42,a44,a46,a48,a50,a52,a54,a56,a58,a60,a62,a64,a66,
a68,a70,a72,a74,a76,a78,a80,a82,a84,a86,a88,a90,a92,a94,a96,
a98,a100,a102,a104,a106,a108,a110,a112,a114,a116,a118,a120,a122,a124,a126,
a128,a130,a132,a134,a136,a138,a140,a142,a144,a146,a148,a150,a152,a154,a156,
a158,a160,a162,a164,a166,a168,a170,a172,a174,a176,a178,a180,a182,a184,a186,
a188,a190,a192,a194,a196,a198,a200,a202,a204,a206,a208,a210,a212,a214,a216,
a218,a220,a222,a224,a226,a228,a230,a232,a234,a236,a238,a240,a242,a244,a246,
a248,a250,a252,a254,a256,a258,a260,a262,a264,a266,a268,a270,a272,a274,a276,
a278,a280,a282,a284,a286,a288,a290,a292,a294,a296,a298,a300,a302,a304,a306,
a308,a310,a312,a314,a316,a318,a320,a322,a324,a326,a328,a330,a332,a334,a336,
a338,a340,a342,a344,a346,a348,a350,a352,a354,a356,a358,a360,a362,a364,a366,
a368,a370,a372,a374,a376,a378,a380,a382,a384,a386,a388,a390,a392,a394,a396,
a398,a400,a402,a404,a406,a408,a410,a412,a414,a416,a418,a420,a422,a424,a426,
a428,a430,a432,a434,a436,a438,a440,a442,a444,a446,a448,a450,a452,a454,a456,
a458,a460,a462,a464,a466,a468,a470,a472,a474,a476,a478,a480,a482,a484,a486,
a488,a490,a492,a494,a496,a498,a500,a502,a504,a506,a508,a510,a512,a514,a516,
a518,a520,a522,a524,a526,a528,a530,a532,a534,a536,a538,a540,a542,a544,a546,
a548,a550,a552,a554,a556,a558,a560,a562,a564,a566,a568,a570,a572,a574,a576,
a578,a580,a582,a584,a586,a588,a590,a592,a594,a596,a598,a600,a602,a604,a606,
a608,a610,a612,a614,a616,a618,a620,a622,a624,a626,a628,a630,a632,a634,a636,
a638,a640,a642,a644,a646,a648,a650,a652,a654,a656,a658,a660,a662,a664,a666,
a668,a670,a672,a674,a676,a678,a680,a682,a684,a686,a688,a690,a692,a694,a696,
a698,a700,a702,a704,a706,a708,a710,a712,a714,a716,a718,a720,a722,a724,a726,
a728,a730,a732,a734,a736,a738,a740,a742,a744,a746,a748,a750,a752,a754,a756,
a758,a760,a762,a764,a766,a768,a770,a772,a774,a776,a778,a780,a782,a784,a786,
a788,a790,a792,a794,a796,a798,a800,a802,a804,a806,a808,a810,a812,a814,a816,
a818,a820,a822,a824,a826,a828,a830,a832,a834,a836,a838,a840,a842,a844,a846,
a848,a850,a852,a854,a856,a858,a860,a862,a864,a866,a868,a870,a872,a874,a876,
a878,a880,a882,a884,a886,a888,a890,a892,a894,a896,a898,a900,a902,a904,a906,
a908,a910,a912,a914,a916,a918,a920,a922,a924,a926,a928,a930,a932,a934,a936,
a938,a940,a942,a944,a946,a948,a950,a952,a954,a956,a958,a960,a962,a964,a966,
a968,a970,a972,a974,a976,a978,a980,a982,a984,a986,a988,a990,a992,a994,a996,
a998,a1000,a1002,a1004,a1006,a1008,a1010,a1012,a1014,a1016,a1018,a1020,a1022,a1024,a1026,
a1028,a1030,a1032,a1034,a1036,a1038,a1040,a1042,a1044,a1046,a1048,a1050,a1052,a1054,a1056,
a1058,a1060,a1062,a1064,a1066,a1068,a1070,a1072,a1074,a1076,a1078,a1080,a1082,a1084,a1086,
a1088,a1090,a1092,a1094,a1096,a1098,a1100,a1102,a1104,a1106,a1108,a1110,a1112,a1114,a1116,
a1118,a1120,a1122,a1124,a1126,a1128,a1130,a1132,a1134,a1136,a1138,a1140,a1142,a1144,a1146,
a1148,a1150,a1152,a1154,a1156,a1158,a1160,a1162,a1164,a1166,a1168,a1170,a1172,a1174,a1176,
a1178,a1180,a1182,a1184,a1186,a1188,a1190,a1192,a1194,a1196,a1198,a1200,a1202,a1204,a1206,
a1208,a1210,a1212,a1214,a1216,a1218,a1220,a1222,a1224,a1226,a1228,a1230,a1232,a1234,a1236,
a1238,a1240,a1242,a1244,a1246,a1248,a1250,a1252,a1254,a1256,a1258,a1260,a1262,a1264,a1266,
a1268,a1270,a1272,a1274,a1276,a1278,a1280,a1282,a1284,a1286,a1288,a1290,a1292,a1294,a1296,
a1298,a1300,a1302,a1304,a1306,a1308,a1310,a1312,a1314,a1316,a1318,a1320,a1322,a1324,a1326,
a1328,a1330,a1332,a1334,a1336,a1338,a1340,a1342,a1344,a1346,a1348,a1350,a1352,a1354,a1356,
a1358,a1360,a1362,a1364,a1366,a1368,a1370,a1372,a1374,a1376,a1378,a1380,a1382,a1384,a1386,
a1388,a1390,a1392,a1394,a1396,a1398,a1400,a1402,a1404,a1406,a1408,a1410,a1412,a1414,a1416,
a1418,a1420,a1422,a1424,p0;

reg l6,l8,l10,l12,l14,l16,l18,l20,l22,l24;

initial
begin
   l6 = 0;
   l8 = 0;
   l10 = 0;
   l12 = 0;
   l14 = 0;
   l16 = 0;
   l18 = 0;
   l20 = 0;
   l22 = 0;
   l24 = 0;
end

always @(posedge na162)
   l6 <= na162;

always @(posedge i2)
   l8 <= i2;

always @(posedge na228)
   l10 <= na228;

always @(posedge na776)
   l12 <= na776;

always @(posedge na800)
   l14 <= na800;

always @(posedge na822)
   l16 <= na822;

always @(posedge na1334)
   l18 <= na1334;

always @(posedge na1358)
   l20 <= na1358;

always @(posedge na1380)
   l22 <= na1380;

always @(posedge na1424)
   l24 <= na1424;


assign na162 = ~a162;
assign na228 = ~a228;
assign na776 = ~a776;
assign na800 = ~a800;
assign na822 = ~a822;
assign na1334 = ~a1334;
assign na1358 = ~a1358;
assign na1380 = ~a1380;
assign na1424 = ~a1424;
assign a26 = ~l20 & l18;
assign a28 = ~a26 & l18;
assign a30 = l14 & ~l12;
assign a32 = ~a30 & l14;
assign a34 = ~a32 & ~a28;
assign a36 = a34 & l16;
assign a38 = ~l14 & l12;
assign a40 = ~a38 & l12;
assign a42 = l20 & ~l18;
assign a44 = ~a42 & l20;
assign a46 = ~a44 & ~a40;
assign a48 = ~a28 & l14;
assign a50 = a48 & ~l12;
assign a52 = ~a28 & l12;
assign a54 = a52 & ~l14;
assign a56 = a54 & ~a50;
assign a58 = a56 & ~a36;
assign a60 = a46 & l22;
assign a62 = a42 & ~l12;
assign a64 = a42 & l12;
assign a66 = a64 & ~l14;
assign a68 = ~a66 & ~a62;
assign a70 = a26 & l12;
assign a72 = a70 & ~l14;
assign a74 = a26 & ~l12;
assign a76 = ~a74 & ~a72;
assign a78 = ~a76 & a68;
assign a80 = a78 & ~a60;
assign a82 = a80 & a58;
assign a84 = a34 & ~i2;
assign a86 = a84 & l16;
assign a88 = a46 & i2;
assign a90 = a88 & l22;
assign a92 = ~a90 & ~a86;
assign a94 = ~a28 & ~i2;
assign a96 = a94 & l14;
assign a98 = ~l18 & i2;
assign a100 = a98 & l20;
assign a102 = ~a100 & ~a96;
assign a104 = ~a102 & ~l12;
assign a106 = a100 & l12;
assign a108 = a106 & ~l14;
assign a110 = ~a108 & ~a104;
assign a112 = l18 & i2;
assign a114 = a112 & ~l20;
assign a116 = ~a114 & ~a94;
assign a118 = ~a116 & l12;
assign a120 = a118 & ~l14;
assign a122 = a114 & ~l12;
assign a124 = ~a122 & ~a120;
assign a126 = a124 & a110;
assign a128 = a124 & ~a110;
assign a130 = a126 & a92;
assign a132 = a126 & ~a92;
assign a134 = a128 & a92;
assign a136 = ~a132 & ~a130;
assign a138 = a136 & a134;
assign a140 = ~a134 & l6;
assign a142 = a134 & ~i2;
assign a144 = ~a142 & ~a140;
assign a146 = ~a144 & ~a132;
assign a148 = a132 & l6;
assign a150 = ~a148 & ~a146;
assign a152 = ~a150 & ~a130;
assign a154 = a130 & l6;
assign a156 = ~a154 & ~a152;
assign a158 = ~a156 & a138;
assign a160 = ~a138 & l6;
assign a162 = ~a160 & ~a158;
assign a164 = a128 & ~a92;
assign a166 = ~a124 & a110;
assign a168 = a166 & a92;
assign a170 = a166 & ~a92;
assign a172 = ~a134 & ~a132;
assign a174 = a170 & ~a168;
assign a176 = a174 & ~a164;
assign a178 = a176 & a172;
assign a180 = ~a178 & ~a132;
assign a182 = ~a180 & ~a130;
assign a184 = l10 & i2;
assign a186 = ~a184 & i2;
assign a188 = ~a170 & l10;
assign a190 = a184 & a170;
assign a192 = ~a190 & ~a188;
assign a194 = ~a192 & ~a168;
assign a196 = a168 & l10;
assign a198 = ~a196 & ~a194;
assign a200 = ~a198 & ~a164;
assign a202 = a164 & l10;
assign a204 = ~a202 & ~a200;
assign a206 = ~a204 & ~a134;
assign a208 = a134 & l10;
assign a210 = ~a208 & ~a206;
assign a212 = ~a210 & ~a132;
assign a214 = ~a186 & a132;
assign a216 = ~a214 & ~a212;
assign a218 = ~a216 & ~a130;
assign a220 = a130 & l10;
assign a222 = ~a220 & ~a218;
assign a224 = ~a222 & a182;
assign a226 = ~a182 & l10;
assign a228 = ~a226 & ~a224;
assign a230 = l24 & ~i2;
assign a232 = ~a230 & ~a184;
assign a234 = ~l6 & i2;
assign a236 = l6 & ~i2;
assign a238 = ~a236 & ~a234;
assign a240 = ~a238 & ~a232;
assign a242 = a130 & ~i4;
assign a244 = a168 & ~i4;
assign a246 = ~a244 & ~a174;
assign a248 = ~a246 & ~a164;
assign a250 = ~a240 & a164;
assign a252 = ~a250 & ~a248;
assign a254 = ~a252 & ~a134;
assign a256 = ~a254 & ~a134;
assign a258 = ~a256 & ~a132;
assign a260 = ~a258 & ~a132;
assign a262 = ~a260 & ~a130;
assign a264 = ~a262 & ~a242;
assign a266 = ~a40 & ~i2;
assign a268 = ~a32 & i2;
assign a270 = a268 & l16;
assign a272 = ~a270 & ~a266;
assign a274 = ~l12 & i2;
assign a276 = a274 & l14;
assign a278 = l12 & i2;
assign a280 = a278 & ~l14;
assign a282 = ~a280 & ~a266;
assign a284 = ~a280 & a276;
assign a286 = ~a284 & a276;
assign a288 = ~a286 & ~a40;
assign a290 = a288 & ~i4;
assign a292 = a290 & ~a272;
assign a294 = a280 & ~a276;
assign a296 = ~a294 & a280;
assign a298 = ~a296 & ~a32;
assign a300 = a298 & i4;
assign a302 = a300 & l16;
assign a304 = ~a302 & ~a292;
assign a306 = ~a40 & ~i4;
assign a308 = a306 & a276;
assign a310 = ~l12 & i4;
assign a312 = a310 & l14;
assign a314 = ~a312 & ~a308;
assign a316 = ~a314 & ~a280;
assign a318 = a312 & a280;
assign a320 = a318 & ~a276;
assign a322 = ~a320 & ~a316;
assign a324 = l12 & i4;
assign a326 = a324 & ~l14;
assign a328 = ~a326 & ~a306;
assign a330 = ~a328 & a280;
assign a332 = a330 & ~a276;
assign a334 = a326 & ~a280;
assign a336 = ~a334 & ~a332;
assign a338 = ~a276 & ~a266;
assign a340 = a282 & a276;
assign a342 = ~a340 & a276;
assign a344 = ~a342 & ~a40;
assign a346 = a344 & ~a240;
assign a348 = a346 & a270;
assign a350 = ~a282 & ~a276;
assign a352 = ~a350 & ~a282;
assign a354 = ~a352 & ~a32;
assign a356 = a354 & a240;
assign a358 = a356 & l16;
assign a360 = ~a358 & ~a348;
assign a362 = ~a240 & ~a40;
assign a364 = a362 & a276;
assign a366 = a240 & ~l12;
assign a368 = a366 & l14;
assign a370 = ~a368 & ~a364;
assign a372 = ~a370 & a282;
assign a374 = a368 & ~a282;
assign a376 = a374 & ~a276;
assign a378 = ~a376 & ~a372;
assign a380 = a240 & l12;
assign a382 = a380 & ~l14;
assign a384 = ~a382 & ~a362;
assign a386 = ~a384 & ~a282;
assign a388 = a386 & ~a276;
assign a390 = a382 & a282;
assign a392 = ~a390 & ~a388;
assign a394 = a344 & ~i4;
assign a396 = a394 & ~a272;
assign a398 = a354 & i4;
assign a400 = a398 & l16;
assign a402 = ~a400 & ~a396;
assign a404 = ~a314 & a282;
assign a406 = a312 & ~a282;
assign a408 = a406 & ~a276;
assign a410 = ~a408 & ~a404;
assign a412 = ~a328 & ~a282;
assign a414 = a412 & ~a276;
assign a416 = a326 & a282;
assign a418 = ~a416 & ~a414;
assign a420 = a288 & a170;
assign a422 = a420 & a270;
assign a424 = a298 & ~a170;
assign a426 = a424 & l16;
assign a428 = ~a426 & ~a422;
assign a430 = a170 & ~a40;
assign a432 = a430 & a276;
assign a434 = ~a170 & ~l12;
assign a436 = a434 & l14;
assign a438 = ~a436 & ~a432;
assign a440 = ~a438 & ~a280;
assign a442 = a436 & a280;
assign a444 = a442 & ~a276;
assign a446 = ~a444 & ~a440;
assign a448 = ~a170 & l12;
assign a450 = a448 & ~l14;
assign a452 = ~a450 & ~a430;
assign a454 = ~a452 & a280;
assign a456 = a454 & ~a276;
assign a458 = a450 & ~a280;
assign a460 = ~a458 & ~a456;
assign a462 = ~a460 & a446;
assign a464 = ~a462 & ~a460;
assign a466 = a418 & ~a410;
assign a468 = ~a466 & ~a410;
assign a470 = ~a468 & ~a464;
assign a472 = a470 & a168;
assign a474 = a472 & ~a402;
assign a476 = ~a418 & a410;
assign a478 = ~a476 & ~a418;
assign a480 = a460 & ~a446;
assign a482 = ~a480 & ~a446;
assign a484 = ~a482 & ~a478;
assign a486 = a484 & ~a168;
assign a488 = a486 & ~a428;
assign a490 = ~a488 & ~a474;
assign a492 = ~a464 & a168;
assign a494 = a492 & ~a410;
assign a496 = a460 & ~a168;
assign a498 = a496 & ~a446;
assign a500 = ~a498 & ~a494;
assign a502 = ~a500 & a418;
assign a504 = a498 & ~a418;
assign a506 = a504 & a410;
assign a508 = ~a506 & ~a502;
assign a510 = ~a460 & ~a168;
assign a512 = a510 & a446;
assign a514 = ~a512 & ~a492;
assign a516 = ~a514 & ~a418;
assign a518 = a516 & a410;
assign a520 = a512 & a418;
assign a522 = ~a520 & ~a518;
assign a524 = ~a522 & a508;
assign a526 = ~a524 & ~a522;
assign a528 = a392 & ~a378;
assign a530 = ~a528 & ~a378;
assign a532 = ~a530 & ~a526;
assign a534 = a532 & a164;
assign a536 = a534 & ~a360;
assign a538 = ~a392 & a378;
assign a540 = ~a538 & ~a392;
assign a542 = a522 & ~a508;
assign a544 = ~a542 & ~a508;
assign a546 = ~a544 & ~a540;
assign a548 = a546 & ~a164;
assign a550 = a548 & ~a490;
assign a552 = ~a550 & ~a536;
assign a554 = ~a526 & a164;
assign a556 = a554 & ~a378;
assign a558 = a522 & ~a164;
assign a560 = a558 & ~a508;
assign a562 = ~a560 & ~a556;
assign a564 = ~a562 & a392;
assign a566 = a560 & ~a392;
assign a568 = a566 & a378;
assign a570 = ~a568 & ~a564;
assign a572 = ~a522 & ~a164;
assign a574 = a572 & a508;
assign a576 = ~a574 & ~a554;
assign a578 = ~a576 & ~a392;
assign a580 = a578 & a378;
assign a582 = a574 & a392;
assign a584 = ~a582 & ~a580;
assign a586 = ~a584 & a570;
assign a588 = ~a586 & ~a584;
assign a590 = ~a338 & ~a280;
assign a592 = ~a590 & ~a338;
assign a594 = ~a592 & ~a588;
assign a596 = a594 & a134;
assign a598 = a596 & ~a272;
assign a600 = a338 & a280;
assign a602 = ~a600 & a280;
assign a604 = a584 & ~a570;
assign a606 = ~a604 & ~a570;
assign a608 = ~a606 & ~a602;
assign a610 = a608 & ~a134;
assign a612 = a610 & ~a552;
assign a614 = ~a612 & ~a598;
assign a616 = ~a588 & a134;
assign a618 = a616 & ~a338;
assign a620 = a584 & ~a134;
assign a622 = a620 & ~a570;
assign a624 = ~a622 & ~a618;
assign a626 = ~a624 & ~a280;
assign a628 = a622 & a280;
assign a630 = a628 & a338;
assign a632 = ~a630 & ~a626;
assign a634 = ~a584 & ~a134;
assign a636 = a634 & a570;
assign a638 = ~a636 & ~a616;
assign a640 = ~a638 & a280;
assign a642 = a640 & a338;
assign a644 = a636 & ~a280;
assign a646 = ~a644 & ~a642;
assign a648 = ~a646 & a632;
assign a650 = ~a648 & ~a646;
assign a652 = ~a650 & ~a592;
assign a654 = a652 & a132;
assign a656 = a654 & a270;
assign a658 = a646 & ~a632;
assign a660 = ~a658 & ~a632;
assign a662 = ~a660 & ~a602;
assign a664 = a662 & ~a132;
assign a666 = a664 & ~a614;
assign a668 = ~a666 & ~a656;
assign a670 = ~a650 & a132;
assign a672 = a670 & ~a338;
assign a674 = a646 & ~a132;
assign a676 = a674 & ~a632;
assign a678 = ~a676 & ~a672;
assign a680 = ~a678 & ~a280;
assign a682 = a676 & a280;
assign a684 = a682 & a338;
assign a686 = ~a684 & ~a680;
assign a688 = ~a646 & ~a132;
assign a690 = a688 & a632;
assign a692 = ~a690 & ~a670;
assign a694 = ~a692 & a280;
assign a696 = a694 & a338;
assign a698 = a690 & ~a280;
assign a700 = ~a698 & ~a696;
assign a702 = ~a700 & a686;
assign a704 = ~a702 & ~a700;
assign a706 = a336 & ~a322;
assign a708 = ~a706 & ~a322;
assign a710 = ~a708 & ~a704;
assign a712 = a710 & a130;
assign a714 = a712 & ~a304;
assign a716 = ~a336 & a322;
assign a718 = ~a716 & ~a336;
assign a720 = a700 & ~a686;
assign a722 = ~a720 & ~a686;
assign a724 = ~a722 & ~a718;
assign a726 = a724 & ~a130;
assign a728 = a726 & ~a668;
assign a730 = ~a728 & ~a714;
assign a732 = ~a704 & a130;
assign a734 = a732 & ~a322;
assign a736 = a700 & ~a130;
assign a738 = a736 & ~a686;
assign a740 = ~a738 & ~a734;
assign a742 = ~a740 & a336;
assign a744 = a738 & ~a336;
assign a746 = a744 & a322;
assign a748 = ~a746 & ~a742;
assign a750 = ~a700 & ~a130;
assign a752 = a750 & a686;
assign a754 = ~a752 & ~a732;
assign a756 = ~a754 & ~a336;
assign a758 = a756 & a322;
assign a760 = a752 & a336;
assign a762 = ~a760 & ~a758;
assign a764 = ~a264 & ~l12;
assign a766 = ~a764 & ~a38;
assign a768 = ~a766 & ~a762;
assign a770 = a768 & a748;
assign a772 = a762 & a38;
assign a774 = a772 & a264;
assign a776 = ~a774 & ~a770;
assign a778 = ~a748 & ~a264;
assign a780 = a264 & l14;
assign a782 = ~a780 & ~a778;
assign a784 = ~a782 & ~l12;
assign a786 = ~a748 & a38;
assign a788 = a786 & ~a264;
assign a790 = ~a788 & ~a784;
assign a792 = ~a790 & a762;
assign a794 = ~a762 & a30;
assign a796 = a794 & a748;
assign a798 = a796 & a264;
assign a800 = ~a798 & ~a792;
assign a802 = a762 & ~a748;
assign a804 = ~a802 & ~a748;
assign a806 = ~a804 & ~a40;
assign a808 = a806 & ~a730;
assign a810 = a808 & ~a264;
assign a812 = ~a762 & a748;
assign a814 = ~a812 & ~a762;
assign a816 = ~a814 & ~a32;
assign a818 = a816 & l16;
assign a820 = a818 & a264;
assign a822 = ~a820 & ~a810;
assign a824 = ~a28 & i2;
assign a826 = ~a44 & ~i2;
assign a828 = a826 & l22;
assign a830 = ~a828 & ~a824;
assign a832 = ~l18 & ~i2;
assign a834 = a832 & l20;
assign a836 = l18 & ~i2;
assign a838 = a836 & ~l20;
assign a840 = ~a838 & ~a824;
assign a842 = ~a838 & a834;
assign a844 = ~a842 & a834;
assign a846 = ~a844 & ~a28;
assign a848 = a846 & ~i4;
assign a850 = a848 & ~a830;
assign a852 = a838 & ~a834;
assign a854 = ~a852 & a838;
assign a856 = ~a854 & ~a44;
assign a858 = a856 & i4;
assign a860 = a858 & l22;
assign a862 = ~a860 & ~a850;
assign a864 = ~a28 & ~i4;
assign a866 = a864 & a834;
assign a868 = ~l18 & i4;
assign a870 = a868 & l20;
assign a872 = ~a870 & ~a866;
assign a874 = ~a872 & ~a838;
assign a876 = a870 & a838;
assign a878 = a876 & ~a834;
assign a880 = ~a878 & ~a874;
assign a882 = l18 & i4;
assign a884 = a882 & ~l20;
assign a886 = ~a884 & ~a864;
assign a888 = ~a886 & a838;
assign a890 = a888 & ~a834;
assign a892 = a884 & ~a838;
assign a894 = ~a892 & ~a890;
assign a896 = ~a834 & ~a824;
assign a898 = a840 & a834;
assign a900 = ~a898 & a834;
assign a902 = ~a900 & ~a28;
assign a904 = a902 & ~a240;
assign a906 = a904 & a828;
assign a908 = ~a840 & ~a834;
assign a910 = ~a908 & ~a840;
assign a912 = ~a910 & ~a44;
assign a914 = a912 & a240;
assign a916 = a914 & l22;
assign a918 = ~a916 & ~a906;
assign a920 = ~a240 & ~a28;
assign a922 = a920 & a834;
assign a924 = a240 & ~l18;
assign a926 = a924 & l20;
assign a928 = ~a926 & ~a922;
assign a930 = ~a928 & a840;
assign a932 = a926 & ~a840;
assign a934 = a932 & ~a834;
assign a936 = ~a934 & ~a930;
assign a938 = a240 & l18;
assign a940 = a938 & ~l20;
assign a942 = ~a940 & ~a920;
assign a944 = ~a942 & ~a840;
assign a946 = a944 & ~a834;
assign a948 = a940 & a840;
assign a950 = ~a948 & ~a946;
assign a952 = a902 & ~i4;
assign a954 = a952 & ~a830;
assign a956 = a912 & i4;
assign a958 = a956 & l22;
assign a960 = ~a958 & ~a954;
assign a962 = ~a872 & a840;
assign a964 = a870 & ~a840;
assign a966 = a964 & ~a834;
assign a968 = ~a966 & ~a962;
assign a970 = ~a886 & ~a840;
assign a972 = a970 & ~a834;
assign a974 = a884 & a840;
assign a976 = ~a974 & ~a972;
assign a978 = a846 & a170;
assign a980 = a978 & a828;
assign a982 = a856 & ~a170;
assign a984 = a982 & l22;
assign a986 = ~a984 & ~a980;
assign a988 = a170 & ~a28;
assign a990 = a988 & a834;
assign a992 = ~a170 & ~l18;
assign a994 = a992 & l20;
assign a996 = ~a994 & ~a990;
assign a998 = ~a996 & ~a838;
assign a1000 = a994 & a838;
assign a1002 = a1000 & ~a834;
assign a1004 = ~a1002 & ~a998;
assign a1006 = ~a170 & l18;
assign a1008 = a1006 & ~l20;
assign a1010 = ~a1008 & ~a988;
assign a1012 = ~a1010 & a838;
assign a1014 = a1012 & ~a834;
assign a1016 = a1008 & ~a838;
assign a1018 = ~a1016 & ~a1014;
assign a1020 = ~a1018 & a1004;
assign a1022 = ~a1020 & ~a1018;
assign a1024 = a976 & ~a968;
assign a1026 = ~a1024 & ~a968;
assign a1028 = ~a1026 & ~a1022;
assign a1030 = a1028 & a168;
assign a1032 = a1030 & ~a960;
assign a1034 = ~a976 & a968;
assign a1036 = ~a1034 & ~a976;
assign a1038 = a1018 & ~a1004;
assign a1040 = ~a1038 & ~a1004;
assign a1042 = ~a1040 & ~a1036;
assign a1044 = a1042 & ~a168;
assign a1046 = a1044 & ~a986;
assign a1048 = ~a1046 & ~a1032;
assign a1050 = ~a1022 & a168;
assign a1052 = a1050 & ~a968;
assign a1054 = a1018 & ~a168;
assign a1056 = a1054 & ~a1004;
assign a1058 = ~a1056 & ~a1052;
assign a1060 = ~a1058 & a976;
assign a1062 = a1056 & ~a976;
assign a1064 = a1062 & a968;
assign a1066 = ~a1064 & ~a1060;
assign a1068 = ~a1018 & ~a168;
assign a1070 = a1068 & a1004;
assign a1072 = ~a1070 & ~a1050;
assign a1074 = ~a1072 & ~a976;
assign a1076 = a1074 & a968;
assign a1078 = a1070 & a976;
assign a1080 = ~a1078 & ~a1076;
assign a1082 = ~a1080 & a1066;
assign a1084 = ~a1082 & ~a1080;
assign a1086 = a950 & ~a936;
assign a1088 = ~a1086 & ~a936;
assign a1090 = ~a1088 & ~a1084;
assign a1092 = a1090 & a164;
assign a1094 = a1092 & ~a918;
assign a1096 = ~a950 & a936;
assign a1098 = ~a1096 & ~a950;
assign a1100 = a1080 & ~a1066;
assign a1102 = ~a1100 & ~a1066;
assign a1104 = ~a1102 & ~a1098;
assign a1106 = a1104 & ~a164;
assign a1108 = a1106 & ~a1048;
assign a1110 = ~a1108 & ~a1094;
assign a1112 = ~a1084 & a164;
assign a1114 = a1112 & ~a936;
assign a1116 = a1080 & ~a164;
assign a1118 = a1116 & ~a1066;
assign a1120 = ~a1118 & ~a1114;
assign a1122 = ~a1120 & a950;
assign a1124 = a1118 & ~a950;
assign a1126 = a1124 & a936;
assign a1128 = ~a1126 & ~a1122;
assign a1130 = ~a1080 & ~a164;
assign a1132 = a1130 & a1066;
assign a1134 = ~a1132 & ~a1112;
assign a1136 = ~a1134 & ~a950;
assign a1138 = a1136 & a936;
assign a1140 = a1132 & a950;
assign a1142 = ~a1140 & ~a1138;
assign a1144 = ~a1142 & a1128;
assign a1146 = ~a1144 & ~a1142;
assign a1148 = ~a896 & ~a838;
assign a1150 = ~a1148 & ~a896;
assign a1152 = ~a1150 & ~a1146;
assign a1154 = a1152 & a134;
assign a1156 = a1154 & ~a830;
assign a1158 = a896 & a838;
assign a1160 = ~a1158 & a838;
assign a1162 = a1142 & ~a1128;
assign a1164 = ~a1162 & ~a1128;
assign a1166 = ~a1164 & ~a1160;
assign a1168 = a1166 & ~a134;
assign a1170 = a1168 & ~a1110;
assign a1172 = ~a1170 & ~a1156;
assign a1174 = ~a1146 & a134;
assign a1176 = a1174 & ~a896;
assign a1178 = a1142 & ~a134;
assign a1180 = a1178 & ~a1128;
assign a1182 = ~a1180 & ~a1176;
assign a1184 = ~a1182 & ~a838;
assign a1186 = a1180 & a838;
assign a1188 = a1186 & a896;
assign a1190 = ~a1188 & ~a1184;
assign a1192 = ~a1142 & ~a134;
assign a1194 = a1192 & a1128;
assign a1196 = ~a1194 & ~a1174;
assign a1198 = ~a1196 & a838;
assign a1200 = a1198 & a896;
assign a1202 = a1194 & ~a838;
assign a1204 = ~a1202 & ~a1200;
assign a1206 = ~a1204 & a1190;
assign a1208 = ~a1206 & ~a1204;
assign a1210 = ~a1208 & ~a1150;
assign a1212 = a1210 & a132;
assign a1214 = a1212 & a828;
assign a1216 = a1204 & ~a1190;
assign a1218 = ~a1216 & ~a1190;
assign a1220 = ~a1218 & ~a1160;
assign a1222 = a1220 & ~a132;
assign a1224 = a1222 & ~a1172;
assign a1226 = ~a1224 & ~a1214;
assign a1228 = ~a1208 & a132;
assign a1230 = a1228 & ~a896;
assign a1232 = a1204 & ~a132;
assign a1234 = a1232 & ~a1190;
assign a1236 = ~a1234 & ~a1230;
assign a1238 = ~a1236 & ~a838;
assign a1240 = a1234 & a838;
assign a1242 = a1240 & a896;
assign a1244 = ~a1242 & ~a1238;
assign a1246 = ~a1204 & ~a132;
assign a1248 = a1246 & a1190;
assign a1250 = ~a1248 & ~a1228;
assign a1252 = ~a1250 & a838;
assign a1254 = a1252 & a896;
assign a1256 = a1248 & ~a838;
assign a1258 = ~a1256 & ~a1254;
assign a1260 = ~a1258 & a1244;
assign a1262 = ~a1260 & ~a1258;
assign a1264 = a894 & ~a880;
assign a1266 = ~a1264 & ~a880;
assign a1268 = ~a1266 & ~a1262;
assign a1270 = a1268 & a130;
assign a1272 = a1270 & ~a862;
assign a1274 = ~a894 & a880;
assign a1276 = ~a1274 & ~a894;
assign a1278 = a1258 & ~a1244;
assign a1280 = ~a1278 & ~a1244;
assign a1282 = ~a1280 & ~a1276;
assign a1284 = a1282 & ~a130;
assign a1286 = a1284 & ~a1226;
assign a1288 = ~a1286 & ~a1272;
assign a1290 = ~a1262 & a130;
assign a1292 = a1290 & ~a880;
assign a1294 = a1258 & ~a130;
assign a1296 = a1294 & ~a1244;
assign a1298 = ~a1296 & ~a1292;
assign a1300 = ~a1298 & a894;
assign a1302 = a1296 & ~a894;
assign a1304 = a1302 & a880;
assign a1306 = ~a1304 & ~a1300;
assign a1308 = ~a1258 & ~a130;
assign a1310 = a1308 & a1244;
assign a1312 = ~a1310 & ~a1290;
assign a1314 = ~a1312 & ~a894;
assign a1316 = a1314 & a880;
assign a1318 = a1310 & a894;
assign a1320 = ~a1318 & ~a1316;
assign a1322 = ~a264 & ~l18;
assign a1324 = ~a1322 & ~a26;
assign a1326 = ~a1324 & ~a1320;
assign a1328 = a1326 & a1306;
assign a1330 = a1320 & a26;
assign a1332 = a1330 & a264;
assign a1334 = ~a1332 & ~a1328;
assign a1336 = ~a1306 & ~a264;
assign a1338 = a264 & l20;
assign a1340 = ~a1338 & ~a1336;
assign a1342 = ~a1340 & ~l18;
assign a1344 = ~a1306 & a26;
assign a1346 = a1344 & ~a264;
assign a1348 = ~a1346 & ~a1342;
assign a1350 = ~a1348 & a1320;
assign a1352 = ~a1320 & a42;
assign a1354 = a1352 & a1306;
assign a1356 = a1354 & a264;
assign a1358 = ~a1356 & ~a1350;
assign a1360 = a1320 & ~a1306;
assign a1362 = ~a1360 & ~a1306;
assign a1364 = ~a1362 & ~a28;
assign a1366 = a1364 & ~a1288;
assign a1368 = a1366 & ~a264;
assign a1370 = ~a1320 & a1306;
assign a1372 = ~a1370 & ~a1320;
assign a1374 = ~a1372 & ~a44;
assign a1376 = a1374 & l22;
assign a1378 = a1376 & a264;
assign a1380 = ~a1378 & ~a1368;
assign a1382 = ~a230 & ~i2;
assign a1384 = ~a170 & l24;
assign a1386 = a230 & a170;
assign a1388 = ~a1386 & ~a1384;
assign a1390 = ~a1388 & ~a168;
assign a1392 = a168 & l24;
assign a1394 = ~a1392 & ~a1390;
assign a1396 = ~a1394 & ~a164;
assign a1398 = a164 & l24;
assign a1400 = ~a1398 & ~a1396;
assign a1402 = ~a1400 & ~a134;
assign a1404 = a134 & l24;
assign a1406 = ~a1404 & ~a1402;
assign a1408 = ~a1406 & ~a132;
assign a1410 = ~a1382 & a132;
assign a1412 = ~a1410 & ~a1408;
assign a1414 = ~a1412 & ~a130;
assign a1416 = a130 & l24;
assign a1418 = ~a1416 & ~a1414;
assign a1420 = ~a1418 & a182;
assign a1422 = ~a182 & l24;
assign a1424 = ~a1422 & ~a1420;
assign p0 = a82;

assert property (~p0);

endmodule
