module viseisenberg (i2,i4,i6,i8,i10,i12,i14,p0);

input i2,i4,i6,i8,i10,i12,i14;

output p0;

wire a252,a360,a434,a500,a686,a880,a966,a1040,a1106,a1292,a1338,a1370,a1402,a1424,a1446,
a1482,c1,a60,a62,a64,a66,a68,a70,a72,a74,a76,a78,a80,a82,a84,
a86,a88,a90,a92,a94,a96,a98,a100,a102,a104,a106,a108,a110,a112,a114,
a116,a118,a120,a122,a124,a126,a128,a130,a132,a134,a136,a138,a140,a142,a144,
a146,a148,a150,a152,a154,a156,a158,a160,a162,a164,a166,a168,a170,a172,a174,
a176,a178,a180,a182,a184,a186,a188,a190,a192,a194,a196,a198,a200,a202,a204,
a206,a208,a210,a212,a214,a216,a218,a220,a222,a224,a226,a228,a230,a232,a234,
a236,a238,a240,a242,a244,a246,a248,a250,a254,a256,a258,a260,a262,a264,a266,
a268,a270,a272,a274,a276,a278,a280,a282,a284,a286,a288,a290,a292,a294,a296,
a298,a300,a302,a304,a306,a308,a310,a312,a314,a316,a318,a320,a322,a324,a326,
a328,a330,a332,a334,a336,a338,a340,a342,a344,a346,a348,a350,a352,a354,a356,
a358,a362,a364,a366,a368,a370,a372,a374,a376,a378,a380,a382,a384,a386,a388,
a390,a392,a394,a396,a398,a400,a402,a404,a406,a408,a410,a412,a414,a416,a418,
a420,a422,a424,a426,a428,a430,a432,a436,a438,a440,a442,a444,a446,a448,a450,
a452,a454,a456,a458,a460,a462,a464,a466,a468,a470,a472,a474,a476,a478,a480,
a482,a484,a486,a488,a490,a492,a494,a496,a498,a502,a504,a506,a508,a510,a512,
a514,a516,a518,a520,a522,a524,a526,a528,a530,a532,a534,a536,a538,a540,a542,
a544,a546,a548,a550,a552,a554,a556,a558,a560,a562,a564,a566,a568,a570,a572,
a574,a576,a578,a580,a582,a584,a586,a588,a590,a592,a594,a596,a598,a600,a602,
a604,a606,a608,a610,a612,a614,a616,a618,a620,a622,a624,a626,a628,a630,a632,
a634,a636,a638,a640,a642,a644,a646,a648,a650,a652,a654,a656,a658,a660,a662,
a664,a666,a668,a670,a672,a674,a676,a678,a680,a682,a684,a688,a690,a692,a694,
a696,a698,a700,a702,a704,a706,a708,a710,a712,a714,a716,a718,a720,a722,a724,
a726,a728,a730,a732,a734,a736,a738,a740,a742,a744,a746,a748,a750,a752,a754,
a756,a758,a760,a762,a764,a766,a768,a770,a772,a774,a776,a778,a780,a782,a784,
a786,a788,a790,a792,a794,a796,a798,a800,a802,a804,a806,a808,a810,a812,a814,
a816,a818,a820,a822,a824,a826,a828,a830,a832,a834,a836,a838,a840,a842,a844,
a846,a848,a850,a852,a854,a856,a858,a860,a862,a864,a866,a868,a870,a872,a874,
a876,a878,a882,a884,a886,a888,a890,a892,a894,a896,a898,a900,a902,a904,a906,
a908,a910,a912,a914,a916,a918,a920,a922,a924,a926,a928,a930,a932,a934,a936,
a938,a940,a942,a944,a946,a948,a950,a952,a954,a956,a958,a960,a962,a964,a968,
a970,a972,a974,a976,a978,a980,a982,a984,a986,a988,a990,a992,a994,a996,a998,
a1000,a1002,a1004,a1006,a1008,a1010,a1012,a1014,a1016,a1018,a1020,a1022,a1024,a1026,a1028,
a1030,a1032,a1034,a1036,a1038,a1042,a1044,a1046,a1048,a1050,a1052,a1054,a1056,a1058,a1060,
a1062,a1064,a1066,a1068,a1070,a1072,a1074,a1076,a1078,a1080,a1082,a1084,a1086,a1088,a1090,
a1092,a1094,a1096,a1098,a1100,a1102,a1104,a1108,a1110,a1112,a1114,a1116,a1118,a1120,a1122,
a1124,a1126,a1128,a1130,a1132,a1134,a1136,a1138,a1140,a1142,a1144,a1146,a1148,a1150,a1152,
a1154,a1156,a1158,a1160,a1162,a1164,a1166,a1168,a1170,a1172,a1174,a1176,a1178,a1180,a1182,
a1184,a1186,a1188,a1190,a1192,a1194,a1196,a1198,a1200,a1202,a1204,a1206,a1208,a1210,a1212,
a1214,a1216,a1218,a1220,a1222,a1224,a1226,a1228,a1230,a1232,a1234,a1236,a1238,a1240,a1242,
a1244,a1246,a1248,a1250,a1252,a1254,a1256,a1258,a1260,a1262,a1264,a1266,a1268,a1270,a1272,
a1274,a1276,a1278,a1280,a1282,a1284,a1286,a1288,a1290,a1294,a1296,a1298,a1300,a1302,a1304,
a1306,a1308,a1310,a1312,a1314,a1316,a1318,a1320,a1322,a1324,a1326,a1328,a1330,a1332,a1334,
a1336,a1340,a1342,a1344,a1346,a1348,a1350,a1352,a1354,a1356,a1358,a1360,a1362,a1364,a1366,
a1368,a1372,a1374,a1376,a1378,a1380,a1382,a1384,a1386,a1388,a1390,a1392,a1394,a1396,a1398,
a1400,a1404,a1406,a1408,a1410,a1412,a1414,a1416,a1418,a1420,a1422,a1426,a1428,a1430,a1432,
a1434,a1436,a1438,a1440,a1442,a1444,a1448,a1450,a1452,a1454,a1456,a1458,a1460,a1462,a1464,
a1466,a1468,a1470,a1472,a1474,a1476,a1478,a1480,a1484,a1486,a1488,a1490,a1492,a1494,a1496,
a1498,p0;

reg l16,l18,l20,l22,l24,l26,l28,l30,l32,l34,l36,l38,l40,l42,l44,
l46,l48,l50,l52,l54,l56,l58;

initial
begin
   l16 = 0;
   l18 = 0;
   l20 = 0;
   l22 = 0;
   l24 = 0;
   l26 = 0;
   l28 = 0;
   l30 = 0;
   l32 = 0;
   l34 = 0;
   l36 = 0;
   l38 = 0;
   l40 = 0;
   l42 = 0;
   l44 = 0;
   l46 = 0;
   l48 = 0;
   l50 = 0;
   l52 = 0;
   l54 = 0;
   l56 = 0;
   l58 = 0;
end

always @(posedge i6)
   l16 <= i6;

always @(posedge i8)
   l18 <= i8;

always @(posedge i10)
   l20 <= i10;

always @(posedge a252)
   l22 <= a252;

always @(posedge a360)
   l24 <= a360;

always @(posedge a434)
   l26 <= a434;

always @(posedge a500)
   l28 <= a500;

always @(posedge a686)
   l30 <= a686;

always @(posedge a880)
   l32 <= a880;

always @(posedge a966)
   l34 <= a966;

always @(posedge a1040)
   l36 <= a1040;

always @(posedge a1106)
   l38 <= a1106;

always @(posedge a1292)
   l40 <= a1292;

always @(posedge a1338)
   l42 <= a1338;

always @(posedge a1370)
   l44 <= a1370;

always @(posedge a1402)
   l46 <= a1402;

always @(posedge a1424)
   l48 <= a1424;

always @(posedge a1446)
   l50 <= a1446;

always @(posedge i12)
   l52 <= i12;

always @(posedge i14)
   l54 <= i14;

always @(posedge a1482)
   l56 <= a1482;

always @(posedge c1)
   l58 <= c1;


assign a252 = a250 & l58;
assign a360 = a358 & l58;
assign a434 = a432 & l58;
assign a500 = a498 & l58;
assign a686 = a684 & l58;
assign a880 = a878 & l58;
assign a966 = a964 & l58;
assign a1040 = a1038 & l58;
assign a1106 = a1104 & l58;
assign a1292 = a1290 & l58;
assign a1338 = a1336 & l58;
assign a1370 = a1368 & l58;
assign a1402 = a1400 & l58;
assign a1424 = a1422 & l58;
assign a1446 = a1444 & l58;
assign a1482 = ~a1480 & ~a1462;
assign c1 = 1;
assign a60 = ~l28 & ~l26;
assign a62 = a60 & ~l24;
assign a64 = a62 & ~l22;
assign a66 = a62 & l22;
assign a68 = a60 & l24;
assign a70 = a68 & ~l22;
assign a72 = a68 & l22;
assign a74 = ~l28 & l26;
assign a76 = a74 & ~l24;
assign a78 = a76 & ~l22;
assign a80 = a76 & l22;
assign a82 = a74 & l24;
assign a84 = a82 & ~l22;
assign a86 = a82 & l22;
assign a88 = l28 & ~l26;
assign a90 = a88 & ~l24;
assign a92 = a90 & ~l22;
assign a94 = a90 & l22;
assign a96 = a88 & l24;
assign a98 = a96 & ~l22;
assign a100 = a96 & l22;
assign a102 = l28 & l26;
assign a104 = a102 & ~l24;
assign a106 = a104 & ~l22;
assign a108 = a104 & l22;
assign a110 = a102 & l24;
assign a112 = ~a110 & ~a108;
assign a114 = a112 & ~a106;
assign a116 = a114 & ~a100;
assign a118 = a116 & ~a98;
assign a120 = a118 & ~a94;
assign a122 = a120 & ~a92;
assign a124 = a122 & ~a86;
assign a126 = a124 & ~a84;
assign a128 = a126 & ~a80;
assign a130 = a128 & ~a78;
assign a132 = a130 & ~a72;
assign a134 = a132 & ~a70;
assign a136 = a134 & ~a66;
assign a138 = a136 & ~a64;
assign a140 = ~a138 & l16;
assign a142 = ~l44 & l30;
assign a144 = a142 & l48;
assign a146 = l44 & l30;
assign a148 = ~a146 & ~l48;
assign a150 = ~a148 & ~a144;
assign a152 = ~l46 & l30;
assign a154 = a152 & l50;
assign a156 = l46 & l30;
assign a158 = ~a156 & ~l50;
assign a160 = ~a158 & ~a154;
assign a162 = ~a160 & ~a150;
assign a164 = a110 & ~l22;
assign a166 = ~l22 & ~i2;
assign a168 = ~a110 & l22;
assign a170 = ~a168 & i2;
assign a172 = ~a170 & ~a166;
assign a174 = ~a172 & ~a164;
assign a176 = a174 & ~a108;
assign a178 = a176 & a162;
assign a180 = ~a174 & ~a108;
assign a182 = ~a180 & ~a162;
assign a184 = ~a182 & ~a178;
assign a186 = ~a184 & ~a106;
assign a188 = a186 & ~a100;
assign a190 = a188 & ~i2;
assign a192 = ~a186 & ~a100;
assign a194 = ~a192 & i2;
assign a196 = ~a194 & ~a190;
assign a198 = ~a196 & ~a98;
assign a200 = ~a198 & ~a94;
assign a202 = ~a200 & ~a92;
assign a204 = ~a202 & ~a86;
assign a206 = ~a204 & ~a84;
assign a208 = ~a206 & ~a80;
assign a210 = a208 & ~a78;
assign a212 = ~a210 & ~a72;
assign a214 = a212 & a162;
assign a216 = a210 & ~a72;
assign a218 = ~a216 & ~a162;
assign a220 = ~a218 & ~a214;
assign a222 = ~a220 & ~a70;
assign a224 = a222 & l30;
assign a226 = a220 & ~a70;
assign a228 = ~a226 & ~l30;
assign a230 = ~a228 & ~a224;
assign a232 = a230 & ~a66;
assign a234 = ~a232 & ~a64;
assign a236 = ~l22 & ~l16;
assign a238 = a236 & ~a234;
assign a240 = l22 & ~l16;
assign a242 = ~a240 & a234;
assign a244 = ~a242 & ~a238;
assign a246 = ~a244 & a140;
assign a248 = ~a140 & ~l22;
assign a250 = ~a248 & ~a246;
assign a254 = ~l44 & l42;
assign a256 = a254 & l48;
assign a258 = l44 & l42;
assign a260 = ~a258 & ~l48;
assign a262 = ~a260 & ~a256;
assign a264 = ~l46 & l42;
assign a266 = a264 & l50;
assign a268 = l46 & l42;
assign a270 = ~a268 & ~l50;
assign a272 = ~a270 & ~a266;
assign a274 = ~a272 & ~a262;
assign a276 = ~a274 & l42;
assign a278 = a110 & l22;
assign a280 = ~a278 & ~l24;
assign a282 = a280 & ~i2;
assign a284 = ~a278 & l24;
assign a286 = ~a284 & i2;
assign a288 = ~a286 & ~a282;
assign a290 = ~a288 & ~a164;
assign a292 = a290 & ~a108;
assign a294 = a292 & ~a162;
assign a296 = ~a290 & ~a108;
assign a298 = ~a296 & a162;
assign a300 = ~a298 & ~a294;
assign a302 = a300 & ~a106;
assign a304 = ~a302 & ~a100;
assign a306 = a304 & ~i2;
assign a308 = a302 & ~a100;
assign a310 = ~a308 & i2;
assign a312 = ~a310 & ~a306;
assign a314 = ~a312 & ~a98;
assign a316 = a314 & ~a94;
assign a318 = a316 & ~a276;
assign a320 = ~a314 & ~a94;
assign a322 = ~a320 & a276;
assign a324 = ~a322 & ~a318;
assign a326 = a324 & ~a92;
assign a328 = a326 & ~a86;
assign a330 = ~a328 & ~a84;
assign a332 = a330 & ~a80;
assign a334 = a332 & ~a78;
assign a336 = ~a334 & ~a72;
assign a338 = ~a336 & ~a70;
assign a340 = a338 & ~a66;
assign a342 = ~a340 & ~a64;
assign a344 = ~l24 & ~l16;
assign a346 = a344 & a342;
assign a348 = l24 & ~l16;
assign a350 = ~a348 & ~a342;
assign a352 = ~a350 & ~a346;
assign a354 = ~a352 & a140;
assign a356 = ~a140 & ~l24;
assign a358 = ~a356 & ~a354;
assign a362 = ~a278 & ~l26;
assign a364 = a362 & ~i2;
assign a366 = ~a278 & l26;
assign a368 = ~a366 & i2;
assign a370 = ~a368 & ~a364;
assign a372 = ~a370 & ~a164;
assign a374 = a372 & ~a108;
assign a376 = a374 & ~a106;
assign a378 = a376 & ~a100;
assign a380 = a378 & i2;
assign a382 = ~a376 & ~a100;
assign a384 = ~a382 & ~i2;
assign a386 = ~a384 & ~a380;
assign a388 = a386 & ~a98;
assign a390 = a388 & ~a94;
assign a392 = a390 & ~a92;
assign a394 = a392 & ~a86;
assign a396 = ~a394 & ~a84;
assign a398 = ~a396 & ~a80;
assign a400 = a398 & ~a78;
assign a402 = ~a400 & ~a72;
assign a404 = a402 & ~a70;
assign a406 = a404 & ~l30;
assign a408 = ~a402 & ~a70;
assign a410 = ~a408 & l30;
assign a412 = ~a410 & ~a406;
assign a414 = a412 & ~a66;
assign a416 = a414 & ~a64;
assign a418 = ~l26 & ~l16;
assign a420 = a418 & a416;
assign a422 = l26 & ~l16;
assign a424 = ~a422 & ~a416;
assign a426 = ~a424 & ~a420;
assign a428 = ~a426 & a140;
assign a430 = ~a140 & ~l26;
assign a432 = ~a430 & ~a428;
assign a436 = ~a278 & ~l28;
assign a438 = a436 & ~i2;
assign a440 = ~a278 & l28;
assign a442 = ~a440 & i2;
assign a444 = ~a442 & ~a438;
assign a446 = ~a444 & ~a164;
assign a448 = a446 & ~a108;
assign a450 = a448 & ~a106;
assign a452 = a450 & ~a100;
assign a454 = a452 & ~a98;
assign a456 = a454 & ~a94;
assign a458 = a456 & ~a276;
assign a460 = ~a454 & ~a94;
assign a462 = ~a460 & a276;
assign a464 = ~a462 & ~a458;
assign a466 = ~a464 & ~a92;
assign a468 = a466 & ~a86;
assign a470 = ~a468 & ~a84;
assign a472 = a470 & ~a80;
assign a474 = a472 & ~a78;
assign a476 = a474 & ~a72;
assign a478 = a476 & ~a70;
assign a480 = a478 & ~a66;
assign a482 = a480 & ~a64;
assign a484 = ~l28 & ~l16;
assign a486 = a484 & a482;
assign a488 = l28 & ~l16;
assign a490 = ~a488 & ~a482;
assign a492 = ~a490 & ~a486;
assign a494 = ~a492 & a140;
assign a496 = ~a140 & ~l28;
assign a498 = ~a496 & ~a494;
assign a502 = a162 & a108;
assign a504 = ~a502 & ~a106;
assign a506 = ~a504 & ~a100;
assign a508 = a506 & ~a98;
assign a510 = a508 & ~a94;
assign a512 = a510 & ~a92;
assign a514 = ~a512 & ~a86;
assign a516 = ~a514 & ~a84;
assign a518 = ~a516 & ~a80;
assign a520 = a518 & ~a78;
assign a522 = ~a520 & ~a72;
assign a524 = a522 & ~a70;
assign a526 = ~a524 & ~a66;
assign a528 = ~a526 & ~a64;
assign a530 = a528 & l16;
assign a532 = ~a162 & ~l30;
assign a534 = a162 & l30;
assign a536 = ~a534 & ~a532;
assign a538 = ~a108 & ~l30;
assign a540 = a538 & a536;
assign a542 = ~a108 & l30;
assign a544 = ~a542 & ~a536;
assign a546 = ~a544 & ~a540;
assign a548 = ~a546 & ~a106;
assign a550 = a548 & ~l42;
assign a552 = a546 & ~a106;
assign a554 = ~a552 & l42;
assign a556 = ~a554 & ~a550;
assign a558 = ~a556 & ~a100;
assign a560 = a558 & l30;
assign a562 = a556 & ~a100;
assign a564 = ~a562 & ~l30;
assign a566 = ~a564 & ~a560;
assign a568 = ~a566 & ~a98;
assign a570 = a568 & l30;
assign a572 = a566 & ~a98;
assign a574 = ~a572 & ~l30;
assign a576 = ~a574 & ~a570;
assign a578 = ~a576 & ~a94;
assign a580 = a578 & l30;
assign a582 = a576 & ~a94;
assign a584 = ~a582 & ~l30;
assign a586 = ~a584 & ~a580;
assign a588 = ~a586 & ~a92;
assign a590 = a588 & l30;
assign a592 = a586 & ~a92;
assign a594 = ~a592 & ~l30;
assign a596 = ~a594 & ~a590;
assign a598 = a596 & ~a86;
assign a600 = ~a598 & ~a84;
assign a602 = a600 & l30;
assign a604 = a598 & ~a84;
assign a606 = ~a604 & ~l30;
assign a608 = ~a606 & ~a602;
assign a610 = ~a608 & ~a80;
assign a612 = a610 & ~l30;
assign a614 = a608 & ~a80;
assign a616 = ~a614 & l30;
assign a618 = ~a616 & ~a612;
assign a620 = ~a618 & ~a78;
assign a622 = a620 & l42;
assign a624 = a618 & ~a78;
assign a626 = ~a624 & ~l42;
assign a628 = ~a626 & ~a622;
assign a630 = ~a628 & ~a72;
assign a632 = a630 & l30;
assign a634 = a628 & ~a72;
assign a636 = ~a634 & ~l30;
assign a638 = ~a636 & ~a632;
assign a640 = ~a638 & ~a70;
assign a642 = a640 & l30;
assign a644 = a638 & ~a70;
assign a646 = ~a644 & ~l30;
assign a648 = ~a646 & ~a642;
assign a650 = ~a648 & ~a66;
assign a652 = a650 & l42;
assign a654 = a648 & ~a66;
assign a656 = ~a654 & ~l42;
assign a658 = ~a656 & ~a652;
assign a660 = ~a658 & ~a64;
assign a662 = a660 & l30;
assign a664 = a658 & ~a64;
assign a666 = ~a664 & ~l30;
assign a668 = ~a666 & ~a662;
assign a670 = ~l30 & ~l16;
assign a672 = a670 & a668;
assign a674 = l30 & ~l16;
assign a676 = ~a674 & ~a668;
assign a678 = ~a676 & ~a672;
assign a680 = ~a678 & a530;
assign a682 = ~a530 & ~l30;
assign a684 = ~a682 & ~a680;
assign a688 = ~l38 & ~l36;
assign a690 = a688 & ~l34;
assign a692 = a690 & ~l32;
assign a694 = a690 & l32;
assign a696 = a688 & l34;
assign a698 = a696 & ~l32;
assign a700 = a696 & l32;
assign a702 = ~l38 & l36;
assign a704 = a702 & ~l34;
assign a706 = a704 & ~l32;
assign a708 = a704 & l32;
assign a710 = a702 & l34;
assign a712 = a710 & ~l32;
assign a714 = a710 & l32;
assign a716 = l38 & ~l36;
assign a718 = a716 & ~l34;
assign a720 = a718 & ~l32;
assign a722 = a718 & l32;
assign a724 = a716 & l34;
assign a726 = a724 & ~l32;
assign a728 = a724 & l32;
assign a730 = l38 & l36;
assign a732 = a730 & ~l34;
assign a734 = a732 & ~l32;
assign a736 = a732 & l32;
assign a738 = a730 & l34;
assign a740 = ~a738 & ~a736;
assign a742 = a740 & ~a734;
assign a744 = a742 & ~a728;
assign a746 = a744 & ~a726;
assign a748 = a746 & ~a722;
assign a750 = a748 & ~a720;
assign a752 = a750 & ~a714;
assign a754 = a752 & ~a712;
assign a756 = a754 & ~a708;
assign a758 = a756 & ~a706;
assign a760 = a758 & ~a700;
assign a762 = a760 & ~a698;
assign a764 = a762 & ~a694;
assign a766 = a764 & ~a692;
assign a768 = ~a766 & ~l16;
assign a770 = ~l44 & l40;
assign a772 = a770 & l48;
assign a774 = l44 & l40;
assign a776 = ~a774 & ~l48;
assign a778 = ~a776 & ~a772;
assign a780 = ~l46 & l40;
assign a782 = a780 & l50;
assign a784 = l46 & l40;
assign a786 = ~a784 & ~l50;
assign a788 = ~a786 & ~a782;
assign a790 = ~a788 & ~a778;
assign a792 = a738 & ~l32;
assign a794 = ~l32 & ~i4;
assign a796 = ~a738 & l32;
assign a798 = ~a796 & i4;
assign a800 = ~a798 & ~a794;
assign a802 = ~a800 & ~a792;
assign a804 = a802 & ~a736;
assign a806 = a804 & a790;
assign a808 = ~a802 & ~a736;
assign a810 = ~a808 & ~a790;
assign a812 = ~a810 & ~a806;
assign a814 = ~a812 & ~a734;
assign a816 = a814 & ~a728;
assign a818 = a816 & ~i4;
assign a820 = ~a814 & ~a728;
assign a822 = ~a820 & i4;
assign a824 = ~a822 & ~a818;
assign a826 = ~a824 & ~a726;
assign a828 = ~a826 & ~a722;
assign a830 = ~a828 & ~a720;
assign a832 = ~a830 & ~a714;
assign a834 = ~a832 & ~a712;
assign a836 = ~a834 & ~a708;
assign a838 = a836 & ~a706;
assign a840 = ~a838 & ~a700;
assign a842 = a840 & a790;
assign a844 = a838 & ~a700;
assign a846 = ~a844 & ~a790;
assign a848 = ~a846 & ~a842;
assign a850 = ~a848 & ~a698;
assign a852 = a850 & ~l40;
assign a854 = a848 & ~a698;
assign a856 = ~a854 & l40;
assign a858 = ~a856 & ~a852;
assign a860 = a858 & ~a694;
assign a862 = ~a860 & ~a692;
assign a864 = ~l32 & l16;
assign a866 = a864 & ~a862;
assign a868 = l32 & l16;
assign a870 = ~a868 & a862;
assign a872 = ~a870 & ~a866;
assign a874 = ~a872 & a768;
assign a876 = ~a768 & ~l32;
assign a878 = ~a876 & ~a874;
assign a882 = ~a274 & ~l42;
assign a884 = a738 & l32;
assign a886 = ~a884 & ~l34;
assign a888 = a886 & ~i4;
assign a890 = ~a884 & l34;
assign a892 = ~a890 & i4;
assign a894 = ~a892 & ~a888;
assign a896 = ~a894 & ~a792;
assign a898 = a896 & ~a736;
assign a900 = a898 & ~a790;
assign a902 = ~a896 & ~a736;
assign a904 = ~a902 & a790;
assign a906 = ~a904 & ~a900;
assign a908 = a906 & ~a734;
assign a910 = ~a908 & ~a728;
assign a912 = a910 & ~i4;
assign a914 = a908 & ~a728;
assign a916 = ~a914 & i4;
assign a918 = ~a916 & ~a912;
assign a920 = ~a918 & ~a726;
assign a922 = a920 & ~a722;
assign a924 = a922 & ~a882;
assign a926 = ~a920 & ~a722;
assign a928 = ~a926 & a882;
assign a930 = ~a928 & ~a924;
assign a932 = a930 & ~a720;
assign a934 = a932 & ~a714;
assign a936 = ~a934 & ~a712;
assign a938 = a936 & ~a708;
assign a940 = a938 & ~a706;
assign a942 = ~a940 & ~a700;
assign a944 = ~a942 & ~a698;
assign a946 = a944 & ~a694;
assign a948 = ~a946 & ~a692;
assign a950 = ~l34 & l16;
assign a952 = a950 & a948;
assign a954 = l34 & l16;
assign a956 = ~a954 & ~a948;
assign a958 = ~a956 & ~a952;
assign a960 = ~a958 & a768;
assign a962 = ~a768 & ~l34;
assign a964 = ~a962 & ~a960;
assign a968 = ~a884 & ~l36;
assign a970 = a968 & ~i4;
assign a972 = ~a884 & l36;
assign a974 = ~a972 & i4;
assign a976 = ~a974 & ~a970;
assign a978 = ~a976 & ~a792;
assign a980 = a978 & ~a736;
assign a982 = a980 & ~a734;
assign a984 = a982 & ~a728;
assign a986 = a984 & i4;
assign a988 = ~a982 & ~a728;
assign a990 = ~a988 & ~i4;
assign a992 = ~a990 & ~a986;
assign a994 = a992 & ~a726;
assign a996 = a994 & ~a722;
assign a998 = a996 & ~a720;
assign a1000 = a998 & ~a714;
assign a1002 = ~a1000 & ~a712;
assign a1004 = ~a1002 & ~a708;
assign a1006 = a1004 & ~a706;
assign a1008 = ~a1006 & ~a700;
assign a1010 = a1008 & ~a698;
assign a1012 = a1010 & l40;
assign a1014 = ~a1008 & ~a698;
assign a1016 = ~a1014 & ~l40;
assign a1018 = ~a1016 & ~a1012;
assign a1020 = a1018 & ~a694;
assign a1022 = a1020 & ~a692;
assign a1024 = ~l36 & l16;
assign a1026 = a1024 & a1022;
assign a1028 = l36 & l16;
assign a1030 = ~a1028 & ~a1022;
assign a1032 = ~a1030 & ~a1026;
assign a1034 = ~a1032 & a768;
assign a1036 = ~a768 & ~l36;
assign a1038 = ~a1036 & ~a1034;
assign a1042 = ~a884 & ~l38;
assign a1044 = a1042 & ~i4;
assign a1046 = ~a884 & l38;
assign a1048 = ~a1046 & i4;
assign a1050 = ~a1048 & ~a1044;
assign a1052 = ~a1050 & ~a792;
assign a1054 = a1052 & ~a736;
assign a1056 = a1054 & ~a734;
assign a1058 = a1056 & ~a728;
assign a1060 = a1058 & ~a726;
assign a1062 = a1060 & ~a722;
assign a1064 = a1062 & ~a882;
assign a1066 = ~a1060 & ~a722;
assign a1068 = ~a1066 & a882;
assign a1070 = ~a1068 & ~a1064;
assign a1072 = ~a1070 & ~a720;
assign a1074 = a1072 & ~a714;
assign a1076 = ~a1074 & ~a712;
assign a1078 = a1076 & ~a708;
assign a1080 = a1078 & ~a706;
assign a1082 = a1080 & ~a700;
assign a1084 = a1082 & ~a698;
assign a1086 = a1084 & ~a694;
assign a1088 = a1086 & ~a692;
assign a1090 = ~l38 & l16;
assign a1092 = a1090 & a1088;
assign a1094 = l38 & l16;
assign a1096 = ~a1094 & ~a1088;
assign a1098 = ~a1096 & ~a1092;
assign a1100 = ~a1098 & a768;
assign a1102 = ~a768 & ~l38;
assign a1104 = ~a1102 & ~a1100;
assign a1108 = a790 & a736;
assign a1110 = ~a1108 & ~a734;
assign a1112 = ~a1110 & ~a728;
assign a1114 = a1112 & ~a726;
assign a1116 = a1114 & ~a722;
assign a1118 = a1116 & ~a720;
assign a1120 = ~a1118 & ~a714;
assign a1122 = ~a1120 & ~a712;
assign a1124 = ~a1122 & ~a708;
assign a1126 = a1124 & ~a706;
assign a1128 = ~a1126 & ~a700;
assign a1130 = a1128 & ~a698;
assign a1132 = ~a1130 & ~a694;
assign a1134 = ~a1132 & ~a692;
assign a1136 = a1134 & ~l16;
assign a1138 = ~a790 & ~l40;
assign a1140 = a790 & l40;
assign a1142 = ~a1140 & ~a1138;
assign a1144 = ~a736 & ~l40;
assign a1146 = a1144 & a1142;
assign a1148 = ~a736 & l40;
assign a1150 = ~a1148 & ~a1142;
assign a1152 = ~a1150 & ~a1146;
assign a1154 = ~a1152 & ~a734;
assign a1156 = a1154 & ~l42;
assign a1158 = a1152 & ~a734;
assign a1160 = ~a1158 & l42;
assign a1162 = ~a1160 & ~a1156;
assign a1164 = ~a1162 & ~a728;
assign a1166 = a1164 & l40;
assign a1168 = a1162 & ~a728;
assign a1170 = ~a1168 & ~l40;
assign a1172 = ~a1170 & ~a1166;
assign a1174 = ~a1172 & ~a726;
assign a1176 = a1174 & l40;
assign a1178 = a1172 & ~a726;
assign a1180 = ~a1178 & ~l40;
assign a1182 = ~a1180 & ~a1176;
assign a1184 = ~a1182 & ~a722;
assign a1186 = a1184 & l40;
assign a1188 = a1182 & ~a722;
assign a1190 = ~a1188 & ~l40;
assign a1192 = ~a1190 & ~a1186;
assign a1194 = ~a1192 & ~a720;
assign a1196 = a1194 & l40;
assign a1198 = a1192 & ~a720;
assign a1200 = ~a1198 & ~l40;
assign a1202 = ~a1200 & ~a1196;
assign a1204 = a1202 & ~a714;
assign a1206 = ~a1204 & ~a712;
assign a1208 = a1206 & l40;
assign a1210 = a1204 & ~a712;
assign a1212 = ~a1210 & ~l40;
assign a1214 = ~a1212 & ~a1208;
assign a1216 = ~a1214 & ~a708;
assign a1218 = a1216 & ~l40;
assign a1220 = a1214 & ~a708;
assign a1222 = ~a1220 & l40;
assign a1224 = ~a1222 & ~a1218;
assign a1226 = ~a1224 & ~a706;
assign a1228 = a1226 & l42;
assign a1230 = a1224 & ~a706;
assign a1232 = ~a1230 & ~l42;
assign a1234 = ~a1232 & ~a1228;
assign a1236 = ~a1234 & ~a700;
assign a1238 = a1236 & l40;
assign a1240 = a1234 & ~a700;
assign a1242 = ~a1240 & ~l40;
assign a1244 = ~a1242 & ~a1238;
assign a1246 = ~a1244 & ~a698;
assign a1248 = a1246 & l40;
assign a1250 = a1244 & ~a698;
assign a1252 = ~a1250 & ~l40;
assign a1254 = ~a1252 & ~a1248;
assign a1256 = ~a1254 & ~a694;
assign a1258 = a1256 & l42;
assign a1260 = a1254 & ~a694;
assign a1262 = ~a1260 & ~l42;
assign a1264 = ~a1262 & ~a1258;
assign a1266 = ~a1264 & ~a692;
assign a1268 = a1266 & l40;
assign a1270 = a1264 & ~a692;
assign a1272 = ~a1270 & ~l40;
assign a1274 = ~a1272 & ~a1268;
assign a1276 = ~l40 & l16;
assign a1278 = a1276 & a1274;
assign a1280 = l40 & l16;
assign a1282 = ~a1280 & ~a1274;
assign a1284 = ~a1282 & ~a1278;
assign a1286 = ~a1284 & a1136;
assign a1288 = ~a1136 & ~l40;
assign a1290 = ~a1288 & ~a1286;
assign a1294 = ~a164 & ~l42;
assign a1296 = a1294 & l30;
assign a1298 = ~a164 & l42;
assign a1300 = ~a1298 & ~l30;
assign a1302 = ~a1300 & ~a1296;
assign a1304 = a1302 & ~a98;
assign a1306 = ~a792 & ~l42;
assign a1308 = a1306 & l40;
assign a1310 = ~a792 & l42;
assign a1312 = ~a1310 & ~l40;
assign a1314 = ~a1312 & ~a1308;
assign a1316 = ~a1314 & ~a726;
assign a1318 = ~l42 & l16;
assign a1320 = a1318 & ~a1316;
assign a1322 = l42 & l16;
assign a1324 = ~a1322 & a1316;
assign a1326 = ~a1324 & ~a1320;
assign a1328 = ~a1326 & ~l16;
assign a1330 = a1328 & a1304;
assign a1332 = a1326 & ~l16;
assign a1334 = ~a1332 & ~a1304;
assign a1336 = ~a1334 & ~a1330;
assign a1340 = ~l44 & l16;
assign a1342 = ~a884 & l44;
assign a1344 = ~a1342 & ~a712;
assign a1346 = ~a1344 & ~a692;
assign a1348 = a1346 & a1340;
assign a1350 = l44 & l16;
assign a1352 = ~a1350 & ~a1346;
assign a1354 = ~a1352 & ~a1348;
assign a1356 = ~a1354 & ~l16;
assign a1358 = a1356 & l44;
assign a1360 = a1354 & ~l16;
assign a1362 = ~a1360 & ~l44;
assign a1364 = ~a1362 & ~a1358;
assign a1366 = ~a1364 & ~l16;
assign a1368 = ~a1366 & ~a1340;
assign a1372 = ~l46 & l16;
assign a1374 = ~a884 & l46;
assign a1376 = ~a1374 & ~a712;
assign a1378 = a1376 & ~a692;
assign a1380 = ~a1378 & a1372;
assign a1382 = l46 & l16;
assign a1384 = ~a1382 & a1378;
assign a1386 = ~a1384 & ~a1380;
assign a1388 = ~a1386 & ~l16;
assign a1390 = a1388 & l46;
assign a1392 = a1386 & ~l16;
assign a1394 = ~a1392 & ~l46;
assign a1396 = ~a1394 & ~a1390;
assign a1398 = ~a1396 & ~l16;
assign a1400 = ~a1398 & ~a1372;
assign a1404 = ~l48 & ~l16;
assign a1406 = ~a278 & l48;
assign a1408 = ~a1406 & ~a84;
assign a1410 = ~a1408 & ~a64;
assign a1412 = a1410 & a1404;
assign a1414 = l48 & ~l16;
assign a1416 = ~a1414 & ~a1410;
assign a1418 = ~a1416 & ~a1412;
assign a1420 = ~a1418 & l16;
assign a1422 = ~a1420 & ~a1404;
assign a1426 = ~l50 & ~l16;
assign a1428 = ~a278 & l50;
assign a1430 = ~a1428 & ~a84;
assign a1432 = a1430 & ~a64;
assign a1434 = ~a1432 & a1426;
assign a1436 = l50 & ~l16;
assign a1438 = ~a1436 & a1432;
assign a1440 = ~a1438 & ~a1434;
assign a1442 = ~a1440 & l16;
assign a1444 = ~a1442 & ~a1426;
assign a1448 = ~i12 & i10;
assign a1450 = i12 & ~i10;
assign a1452 = ~a1450 & ~a1448;
assign a1454 = ~i14 & i8;
assign a1456 = i14 & ~i8;
assign a1458 = ~a1456 & ~a1454;
assign a1460 = a1458 & a1452;
assign a1462 = ~a1460 & ~l58;
assign a1464 = ~l16 & ~i12;
assign a1466 = l16 & i12;
assign a1468 = ~a1466 & ~a1464;
assign a1470 = l16 & ~i14;
assign a1472 = ~l16 & i14;
assign a1474 = ~a1472 & ~a1470;
assign a1476 = a1474 & a1468;
assign a1478 = a1476 & l56;
assign a1480 = ~a1478 & l58;
assign a1484 = l24 & l22;
assign a1486 = a1484 & ~l26;
assign a1488 = a1486 & l28;
assign a1490 = l34 & l32;
assign a1492 = a1490 & ~l36;
assign a1494 = a1492 & l38;
assign a1496 = a1494 & a1488;
assign a1498 = a1496 & l56;
assign p0 = a1498;

assert property (~p0);

endmodule
