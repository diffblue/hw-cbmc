// 1800 2017 3.14.2.2
timeunit 100ps / 10fs;
timeprecision 10fs;

module main;
endmodule
