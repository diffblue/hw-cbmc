`define something foobar
`something``_else
